VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;
CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS ON ;


LAYER Metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  MINWIDTH 0.05 ;
  AREA 0.0115 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0    0.05 
    WIDTH 0.1  0.06 
    WIDTH 0.35 0.10 
    WIDTH 0.47 0.13 
    WIDTH 0.63 0.15 ;
  SPACING 0.07 ENDOFLINE 0.07 WITHIN 0.025 ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  MINWIDTH 0.05 ;
  WIDTH 0.05 ;
  AREA 0.014 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0    0.05 
    WIDTH 0.09 0.06 
    WIDTH 0.16 0.10 
    WIDTH 0.47 0.13 
    WIDTH 0.63 0.15 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  MINWIDTH 0.05 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0    0.05 
    WIDTH 0.09 0.06 
    WIDTH 0.16 0.10 
    WIDTH 0.47 0.13 
    WIDTH 0.63 0.15 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  MINWIDTH 0.05 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0    0.05 
    WIDTH 0.09 0.06 
    WIDTH 0.16 0.10 
    WIDTH 0.47 0.13 
    WIDTH 0.63 0.15 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  MINWIDTH 0.05 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0    0.05 
    WIDTH 0.09 0.06 
    WIDTH 0.16 0.10 
    WIDTH 0.47 0.13 
    WIDTH 0.63 0.15 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  MINWIDTH 0.05 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0    0.05 
    WIDTH 0.09 0.06 
    WIDTH 0.16 0.10 
    WIDTH 0.47 0.13 
    WIDTH 0.63 0.15 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.10 ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  MINWIDTH 0.05 ;
  PITCH 0.20 0.20 ;
  WIDTH 0.10 ;
  MINWIDTH 0.10 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.10 
    WIDTH 0.2   0.12
    WIDTH 0.4   0.16
    WIDTH 1.5   0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.10 ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  MINWIDTH 0.46 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.10 
    WIDTH 0.2   0.12
    WIDTH 0.4   0.16
    WIDTH 1.5   0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.46 ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.00 1.00 ;
  WIDTH 0.50 ;
  MINWIDTH 0.46 ;
  AREA 1.00 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.50 
    WIDTH 1.5   0.65
    WIDTH 4.5   1.50
    WIDTH 1.5   0.45 ;
END Metal9

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1C DEFAULT 
    LAYER Metal1 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER Metal1 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA12_1C_V

VIA VIA23_1C DEFAULT 
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C_V

VIA VIA23_1ST_N DEFAULT 
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.325000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA23_1ST_N

VIA VIA23_1ST_S DEFAULT 
    LAYER Metal2 ;
        RECT -0.025000 -0.325000 0.025000 0.055000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA23_1ST_S

VIA VIA34_1C DEFAULT 
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA34_1C_V

VIA VIA34_1ST_E DEFAULT 
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.325000 0.025000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA34_1ST_E

VIA VIA34_1ST_W DEFAULT 
    LAYER Metal3 ;
        RECT -0.325000 -0.025000 0.055000 0.025000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA34_1ST_W

VIA VIA45_1C DEFAULT 
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA45_1C

VIA VIA45_1C_H DEFAULT 
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA45_1C_H

VIA VIA45_1C_V DEFAULT 
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA45_1C_V

VIA VIA45_1ST_N DEFAULT 
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.325000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA45_1ST_N

VIA VIA45_1ST_S DEFAULT 
    LAYER Metal4 ;
        RECT -0.025000 -0.325000 0.025000 0.055000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA45_1ST_S

VIA VIA5_0_VH DEFAULT 
    LAYER Metal5 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via5 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA5_0_VH

VIA VIA6_0_HV DEFAULT 
    LAYER Metal6 ;
        RECT -0.260000 -0.100000 0.260000 0.100000 ;
    LAYER Via6 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal7 ;
        RECT -0.100000 -0.260000 0.100000 0.260000 ;
END VIA6_0_HV

VIA VIA7_0_VH DEFAULT 
    LAYER Metal7 ;
        RECT -0.100000 -0.260000 0.100000 0.260000 ;
    LAYER Via7 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal8 ;
        RECT -0.260000 -0.100000 0.260000 0.100000 ;
END VIA7_0_VH

VIA VIA8_0_VH DEFAULT 
    LAYER Metal8 ;
        RECT -0.250000 -0.260000 0.250000 0.260000 ;
    LAYER Via8 ;
        RECT -0.230000 -0.230000 0.230000 0.230000 ;
    LAYER Metal9 ;
        RECT -0.300000 -0.250000 0.300000 0.250000 ;
END VIA8_0_VH


SITE CoreSite
  CLASS CORE ;
  SIZE 0.135 BY 1.2 ;
END CoreSite


MACRO BUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX16 0 0 ;
  SIZE 3.78 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT  0.14 0.42 1.34 0.47 ;
        RECT  0.14 0.62 0.36 0.68 ;
        RECT  0.14 0.42 0.20 0.68 ;
        RECT  1.29 0.42 1.34 0.57 ;
        END
  END A
  PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT  1.46 0.32 3.67 0.46 ;
        RECT  1.46 0.74 3.67 0.89 ;
        RECT  1.46 0.74 1.51 0.96 ;
        RECT  1.46 0.14 1.51 0.46 ;
        RECT  3.54 0.14 3.67 0.96 ;
        END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.78 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.78 0.06 ;
    END
  END VSS
  OBS
        LAYER Metal1 ;
        RECT  0.03 0.30 1.24 0.35 ;
        RECT  0.03 0.30 0.07 0.81 ;
        RECT  0.03 0.75 1.24 0.81 ;
        RECT  1.19 0.14 1.24 0.35 ;
	RECT  1.19 0.68 1.24 0.81 ;
        RECT  1.49 0.62 3.46 0.68 ;
  END
END BUFX16

MACRO BUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
	PORT
        LAYER Metal1 ;
        RECT  0.17 0.33 0.34 0.40 ;
        RECT  0.17 0.33 0.23 0.62 ;
        END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 0.54 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 0.54 0.06 ;
    END
  END VSS
  PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT  0.37 0.20 0.50 0.28 ;
        RECT  0.45 0.20 0.50 1.04 ;
        RECT  0.23 0.85 0.50 0.91 ;
        RECT  0.23 0.85 0.28 1.04 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT  0.04 0.14 0.17 0.23 ;
        RECT  0.04 0.72 0.36 0.78 ;
        RECT  0.04 0.14 0.09 1.04 ;
        RECT  0.31 0.49 0.36 0.78 ;
    END
END BUFX2

MACRO BUFX8
    CLASS CORE ;
    FOREIGN BUFX8 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.89 BY 1.2 ;
    SYMMETRY X Y ;
  SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT  0.14 0.42 0.53 0.47 ;
        RECT  0.14 0.62 0.36 0.68 ;
        RECT  0.14 0.42 0.20 0.68 ;
        RECT  0.48 0.42 0.53 0.57 ;
        END
    END A
    PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.89 1.2 ;
    END
  END VDD

    PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.89 0.06 ;
    END
  END VSS

    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT  0.65 0.33 1.85 0.38 ;
        RECT  0.65 0.82 1.85 0.88 ;
        RECT  0.65 0.82 0.70 0.96 ;
        RECT  0.65 0.14 0.70 0.38 ;
        RECT  1.79 0.14 1.85 0.96 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT  0.04 0.30 0.45 0.35 ;
        RECT  0.04 0.30 0.09 0.88 ;
        RECT  0.04 0.82 0.56 0.88 ;
        RECT  0.52 0.68 0.56 0.88 ;
        RECT  0.36 0.14 0.45 0.35 ;
        RECT  0.52 0.68 1.72 0.72 ;
        RECT  1.65 0.51 1.72 0.72 ;
    END
END BUFX8

MACRO INVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
	PORT
        LAYER Metal1 ;
        RECT  0.17 0.40 0.23 0.76 ;
        END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 0.405 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 0.405 0.06 ;
    END
  END VSS
  PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT  0.23 0.14 0.30 0.28 ;
        RECT  0.31 0.23 0.36 0.92 ;
        RECT  0.23 0.23 0.36 0.28 ;
        RECT  0.24 0.86 0.36 0.92 ;
        RECT  0.24 0.86 0.29 1.05 ;
        END
  END Y
END INVX2

MACRO MX2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X2 0 0 ;
  SIZE 1.89 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.47 0.17 1.52 0.28 ;
        RECT 1.50 0.23 1.56 0.91 ;
        RECT 1.50 0.40 1.74 0.46 ;
        RECT 1.66 0.40 1.74 0.53 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.22 0.41 1.30 0.92 ;
        RECT 1.22 0.41 1.40 0.49 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.43 0.54 0.83 ;
        RECT 0.44 0.76 0.62 0.83 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.78 0.34 1.01 ;
        RECT 0.72 0.73 0.80 1.01 ;
        RECT 0.26 0.94 0.80 1.01 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.89 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.89 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.00 0.21 1.10 0.92 ;
        RECT 0.12 0.21 1.10 0.27 ;
        RECT 0.12 0.21 0.17 0.67 ;
  END
END MX2X2

MACRO OAI2BB1X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X2 0 0 ;
  SIZE 1.89 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.15 0.23 0.77 ;
        RECT 0.06 0.48 0.23 0.77 ;
        RECT 0.39 0.71 0.45 0.98 ;
        RECT 0.17 0.15 0.66 0.22 ;
        RECT 0.06 0.71 0.86 0.77 ;
        RECT 0.80 0.71 0.86 0.98 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.37 0.54 0.52 ;
        RECT 0.33 0.37 0.92 0.45 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.02 0.22 1.17 0.30 ;
        RECT 1.08 0.22 1.17 0.45 ;
        RECT 1.08 0.37 1.38 0.45 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.63 0.33 1.72 0.90 ;
        RECT 1.40 0.85 1.72 0.90 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.89 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.89 0.06 ;
    END
  END VSS
END OAI2BB1X2

MACRO ADDFHX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX2 0 0 ;
  SIZE 4.86 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.39 0.72 4.45 0.99 ;
        RECT 4.43 0.24 4.49 0.78 ;
        RECT 4.43 0.30 4.54 0.43 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.30 0.34 0.43 ;
        RECT 0.28 0.24 0.34 0.99 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.36 0.65 1.89 0.71 ;
        RECT 1.83 0.70 1.96 0.88 ;
        RECT 2.93 0.62 2.99 0.76 ;
        RECT 1.83 0.70 2.99 0.76 ;
        RECT 2.93 0.62 3.97 0.68 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.14 0.50 1.26 0.56 ;
        RECT 1.23 0.49 2.46 0.55 ;
        RECT 2.77 0.46 2.83 0.60 ;
        RECT 2.40 0.54 2.83 0.60 ;
        RECT 3.83 0.42 3.96 0.52 ;
        RECT 2.77 0.46 4.13 0.52 ;
        RECT 4.07 0.46 4.13 0.58 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.83 0.23 1.96 0.38 ;
        RECT 1.83 0.32 2.65 0.38 ;
        RECT 2.59 0.40 2.65 0.44 ;
        RECT 2.59 0.40 3.67 0.36 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.86 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.86 0.06 ;
    END
  END VSS
END ADDFHX2

MACRO ADDFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX2 0 0 ;
  SIZE 4.59 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.25 0.32 4.32 0.99 ;
        RECT 4.25 0.40 4.34 0.53 ;
        RECT 4.22 0.83 4.34 0.99 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 0.49 0.24 0.62 ;
        RECT 0.16 0.49 0.44 0.55 ;
        RECT 0.38 0.24 0.44 1.01 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.19 0.61 1.47 0.67 ;
        RECT 2.06 0.62 2.14 0.91 ;
        RECT 1.43 0.62 3.73 0.68 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.97 0.49 1.09 0.54 ;
        RECT 1.03 0.45 1.57 0.51 ;
        RECT 1.53 0.46 3.96 0.52 ;
        RECT 3.83 0.46 3.96 0.70 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 0.23 1.77 0.36 ;
        RECT 1.64 0.30 3.52 0.36 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.59 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.59 0.06 ;
    END
  END VSS
END ADDFX2


MACRO NAND4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X2 0 0 ;
  SIZE 2.430 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.25 1.23 0.31 ;
        RECT 1.19 0.27 2.12 0.33 ;
        RECT 2.06 0.27 2.12 1.00 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.62 0.32 0.99 ;
        RECT 1.86 0.62 1.94 0.99 ;
        RECT 0.26 0.92 1.94 0.99 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 0.63 0.54 0.70 ;
        RECT 0.46 0.59 0.54 0.72 ;
        RECT 0.48 0.59 0.54 0.82 ;
        RECT 1.60 0.64 1.66 0.82 ;
        RECT 0.48 0.76 1.66 0.82 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.42 1.40 0.50 ;
        RECT 1.33 0.42 1.40 0.66 ;
        RECT 0.69 0.61 1.40 0.66 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.42 1.14 0.50 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.430 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.430 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.12 0.21 0.18 0.92 ;
  END

END NAND4X2


MACRO AOI22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X2 0 0 ;
  SIZE 2.565 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.17 0.21 1.23 0.70 ;
        RECT 1.03 0.61 1.23 0.70 ;
        RECT 1.03 0.63 1.49 0.70 ;
        RECT 1.43 0.63 1.49 0.98 ;
        RECT 0.71 0.21 1.69 0.27 ;
        RECT 1.84 0.79 1.90 0.98 ;
        RECT 1.43 0.92 1.90 0.98 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.56 0.74 0.86 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.54 1.74 0.83 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.50 0.38 1.56 0.51 ;
        RECT 1.32 0.46 1.56 0.51 ;
        RECT 1.50 0.38 1.96 0.44 ;
        RECT 1.84 0.38 1.96 0.70 ;
        RECT 1.84 0.61 2.17 0.70 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.42 0.56 0.50 ;
        RECT 0.48 0.37 0.92 0.46 ;
        RECT 0.84 0.44 1.06 0.51 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.565 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.565 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.10 0.21 0.16 0.92 ;
        RECT 0.10 0.60 0.56 0.66 ;
        RECT 0.50 0.60 0.56 0.96 ;
        RECT 0.10 0.21 0.56 0.27 ;
        RECT 1.84 0.21 2.36 0.27 ;
        RECT 2.30 0.21 2.36 0.97 ;
  END
END AOI22X2

MACRO AND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X2 0 0 ;
  SIZE 1.350 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.25 0.92 0.94 ;
        RECT 0.86 0.40 0.94 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.29 0.59 0.72 ;
        RECT 0.51 0.29 0.59 0.94 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 0.55 0.22 0.92 ;
        RECT 0.22 0.29 0.30 0.91 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.350 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.350 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.06 0.25 1.12 0.94 ;
  END
END AND2X2

MACRO AND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X6 0 0 ;
  SIZE 2.430 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.08 0.28 1.14 0.58 ;
        RECT 1.49 0.28 1.55 0.58 ;
        RECT 1.66 0.53 1.72 0.96 ;
        RECT 1.66 0.79 1.74 0.96 ;
        RECT 1.09 0.90 1.98 0.96 ;
        RECT 1.90 0.28 1.96 0.58 ;
        RECT 1.08 0.53 1.96 0.58 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.79 0.56 0.99 ;
        RECT 0.28 0.79 0.66 0.86 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.62 0.18 0.71 ;
        RECT 0.12 0.32 0.18 0.78 ;
        RECT 0.06 0.62 0.82 0.69 ;
        RECT 0.76 0.32 0.82 0.76 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.430 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.430 0.06 ;
    END
  END VSS

END AND2X6

MACRO AND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X4 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.97 0.690 1.03 0.980 ;
        RECT 0.94 0.220 1.06 0.280 ;
        RECT 1.01 0.240 1.52 0.300 ;
        RECT 1.40 0.180 1.46 0.300 ;
        RECT 1.40 0.690 1.46 0.980 ;
        RECT 1.46 0.240 1.52 0.750 ;
        RECT 0.97 0.690 1.52 0.750 ;
        RECT 1.46 0.400 1.54 0.530 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.360 0.74 0.960 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.10 0.300 0.16 0.630 ;
        RECT 0.10 0.420 0.40 0.500 ;
        RECT 0.32 0.420 0.40 0.810 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS

END AND2X4

MACRO AND3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X2 0 0 ;
  SIZE 1.755 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.15 0.280 1.21 0.460 ;
        RECT 1.15 0.400 1.34 0.460 ;
        RECT 1.26 0.400 1.32 0.980 ;
        RECT 1.26 0.400 1.34 0.530 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.83 0.400 0.92 0.960 ;
        RECT 0.83 0.400 0.96 0.480 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.360 0.34 0.630 ;
        RECT 0.26 0.360 0.57 0.440 ;
        RECT 0.49 0.360 0.57 0.630 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.360 0.16 0.840 ;
        RECT 0.06 0.590 0.16 0.840 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.755 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.755 0.06 ;
    END
  END VSS
END AND3X2

MACRO AND3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X4 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.90 0.270 1.01 0.330 ;
        RECT 1.04 0.780 1.10 0.970 ;
        RECT 1.33 0.270 1.52 0.350 ;
        RECT 0.96 0.290 1.52 0.350 ;
        RECT 1.45 0.780 1.51 0.970 ;
        RECT 1.47 0.270 1.52 0.840 ;
        RECT 1.04 0.780 1.52 0.840 ;
        RECT 1.47 0.490 1.74 0.620 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.70 0.510 0.78 0.860 ;
        RECT 0.70 0.780 0.94 0.860 ;
        RECT 0.86 0.780 0.94 0.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.400 0.34 0.530 ;
        RECT 0.26 0.450 0.44 0.530 ;
        RECT 0.36 0.450 0.44 0.800 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.390 0.14 0.890 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS
END AND3X4

MACRO AND4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X2 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.30 0.610 1.36 0.980 ;
        RECT 0.60 0.150 1.46 0.210 ;
        RECT 1.40 0.150 1.46 0.680 ;
        RECT 1.30 0.610 1.46 0.680 ;
        RECT 1.40 0.400 1.54 0.530 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.00 0.480 1.08 0.720 ;
        RECT 1.06 0.580 1.14 0.910 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.400 0.74 0.900 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.410 0.54 0.910 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 0.420 0.36 0.790 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.66 0.25 1.72 0.94 ;
  END
END AND4X2

MACRO AND4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X4 0 0 ;
  SIZE 2.430 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.18 0.280 1.29 0.340 ;
        RECT 1.29 0.790 1.35 0.980 ;
        RECT 1.29 0.790 1.81 0.850 ;
        RECT 1.61 0.280 1.81 0.360 ;
        RECT 1.25 0.300 1.81 0.360 ;
        RECT 1.75 0.280 1.81 0.980 ;
        RECT 1.70 0.790 1.81 0.980 ;
        RECT 1.75 0.400 1.94 0.530 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.00 0.520 1.08 0.760 ;
        RECT 1.06 0.680 1.14 0.960 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.300 0.74 0.800 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.320 0.56 0.540 ;
        RECT 0.48 0.320 0.56 0.800 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.400 0.34 0.790 ;
        RECT 0.28 0.310 0.36 0.530 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.430 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.430 0.06 ;
    END
  END VSS
END AND4X4

MACRO AO21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X2 0 0 ;
  SIZE 1.755 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.20 0.200 1.26 0.460 ;
        RECT 1.26 0.400 1.34 0.530 ;
        RECT 1.27 0.400 1.34 0.980 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.390 0.34 0.890 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.210 0.54 0.340 ;
        RECT 0.54 0.260 0.61 0.630 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.82 0.440 0.94 0.800 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.755 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.755 0.06 ;
    END
  END VSS
END AO21X2

MACRO AO21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X4 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.02 0.170 1.08 0.310 ;
        RECT 1.23 0.650 1.28 0.980 ;
        RECT 1.43 0.170 1.49 0.310 ;
        RECT 1.02 0.250 1.72 0.310 ;
        RECT 1.23 0.650 1.72 0.710 ;
        RECT 1.64 0.810 1.69 0.980 ;
        RECT 1.66 0.250 1.72 0.860 ;
        RECT 1.66 0.400 1.94 0.460 ;
        RECT 1.86 0.400 1.94 0.530 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.390 0.34 0.890 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.410 0.56 0.890 ;
        RECT 0.46 0.590 0.56 0.890 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 0.410 0.76 0.890 ;
        RECT 0.66 0.590 0.76 0.890 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS
END AO21X4

MACRO AO22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X2 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.210 1.52 0.910 ;
        RECT 1.47 0.780 1.54 0.980 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.02 0.460 1.10 0.920 ;
        RECT 1.02 0.750 1.14 0.920 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.430 0.16 0.910 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.400 0.77 0.500 ;
        RECT 0.69 0.400 0.77 0.850 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.590 0.34 0.720 ;
        RECT 0.26 0.610 0.54 0.700 ;
        RECT 0.46 0.610 0.54 0.870 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS
END AO22X2

MACRO AOI2BB1X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X2 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.400 0.14 0.530 ;
        RECT 0.08 0.250 0.14 0.900 ;
        RECT 0.43 0.170 0.49 0.310 ;
        RECT 0.08 0.840 0.69 0.900 ;
        RECT 0.64 0.840 0.69 0.980 ;
        RECT 0.84 0.170 0.90 0.310 ;
        RECT 0.08 0.250 0.90 0.310 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.500 0.54 0.720 ;
        RECT 0.36 0.500 0.96 0.590 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.250 1.14 0.530 ;
        RECT 1.12 0.400 1.20 0.690 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.360 1.54 0.860 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS
END AOI2BB1X2

MACRO AOI2BB1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X4 0 0 ;
  SIZE 2.565 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.270 0.23 0.850 ;
        RECT 0.23 0.800 0.36 0.870 ;
        RECT 0.41 0.190 0.47 0.330 ;
        RECT 0.61 0.800 0.67 0.980 ;
        RECT 0.81 0.190 0.88 0.330 ;
        RECT 0.17 0.800 1.29 0.850 ;
        RECT 1.23 0.190 1.28 0.330 ;
        RECT 1.23 0.800 1.29 0.980 ;
        RECT 1.64 0.190 1.69 0.330 ;
        RECT 0.17 0.270 1.69 0.330 ;
    END
  END Y
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.230 1.94 0.740 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.300 2.34 0.800 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.540 0.54 0.670 ;
        RECT 0.34 0.540 1.75 0.590 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.565 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.565 0.06 ;
    END
  END VSS
END AOI2BB1X4

MACRO AOI31X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X2 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.70 0.240 1.54 0.300 ;
        RECT 1.46 0.500 1.54 0.630 ;
        RECT 1.48 0.240 1.54 0.900 ;
        RECT 1.50 0.840 1.56 0.960 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.71 0.710 1.05 0.840 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.560 0.54 0.820 ;
        RECT 0.38 0.560 1.05 0.610 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.21 0.390 0.28 0.590 ;
        RECT 0.21 0.390 1.22 0.460 ;
        RECT 1.16 0.390 1.22 0.630 ;
        RECT 1.16 0.500 1.34 0.630 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.390 1.94 0.890 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS
END AOI31X2

MACRO BUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX12 0 0 ;
  SIZE 3.240 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.270 0.29 0.840 ;
        RECT 0.26 0.780 0.34 0.980 ;
        RECT 0.69 0.780 0.75 0.980 ;
        RECT 1.10 0.780 1.16 0.980 ;
        RECT 1.51 0.780 1.57 0.980 ;
        RECT 0.23 0.780 1.98 0.840 ;
        RECT 0.23 0.270 1.98 0.340 ;
        RECT 1.92 0.780 1.98 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.600 2.34 1.030 ;
        RECT 2.26 0.600 2.41 0.680 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.240 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.240 0.06 ;
    END
  END VSS

END BUFX12

MACRO BUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX3 0 0 ;
  SIZE 1.350 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.280 0.23 0.420 ;
        RECT 0.21 0.850 0.28 0.980 ;
        RECT 0.26 0.360 0.32 0.910 ;
        RECT 0.26 0.780 0.34 0.910 ;
        RECT 0.54 0.210 0.60 0.420 ;
        RECT 0.17 0.360 0.60 0.420 ;
        RECT 0.21 0.850 0.69 0.910 ;
        RECT 0.58 0.140 0.65 0.270 ;
        RECT 0.62 0.850 0.69 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.520 0.94 1.020 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.350 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.350 0.06 ;
    END
  END VSS

END BUFX3

MACRO INVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX8 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.48 0.320 1.56 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.320 0.25 0.970 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS

END INVX8

MACRO INVX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX3 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.67 0.320 0.74 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.320 0.27 0.980 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 0.945 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 0.945 0.06 ;
    END
  END VSS

END INVX3

MACRO INVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX4 0 0 ;
  SIZE 1.215 BY 1.2 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.87 0.330 0.95 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.320 0.25 0.980 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.215 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.215 0.06 ;
    END
  END VSS
END INVX4


MACRO INVX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX6 0 0 ;
  SIZE 1.350 BY 1.2 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.07 0.300 1.16 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.320 0.25 0.980 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.350 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.350 0.06 ;
    END
  END VSS
END INVX6

MACRO MX2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X6 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.61 0.190 1.67 0.310 ;
        RECT 1.64 0.630 1.69 0.980 ;
        RECT 1.66 0.200 1.71 0.680 ;
        RECT 1.66 0.400 1.74 0.680 ;
        RECT 2.02 0.200 2.08 0.460 ;
        RECT 2.04 0.400 2.10 0.980 ;
        RECT 1.66 0.400 2.47 0.460 ;
        RECT 2.41 0.280 2.47 0.780 ;
        RECT 2.43 0.200 2.49 0.350 ;
        RECT 2.46 0.730 2.52 0.980 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.480 1.34 0.980 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.410 0.66 0.790 ;
        RECT 0.46 0.590 0.66 0.790 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.720 0.36 0.910 ;
        RECT 0.76 0.720 0.84 0.980 ;
        RECT 0.28 0.890 0.84 0.980 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.835 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.835 0.06 ;
    END
  END VSS
END MX2X6

MACRO MX3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X2 0 0 ;
  SIZE 3.375 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.420 0.37 0.500 ;
        RECT 0.31 0.260 0.37 0.750 ;
        RECT 0.35 0.200 0.41 0.320 ;
        RECT 0.35 0.690 0.41 0.980 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.41 0.820 2.48 0.960 ;
        RECT 2.86 0.780 2.94 0.960 ;
        RECT 2.41 0.870 2.94 0.960 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.40 0.540 2.74 0.620 ;
        RECT 2.66 0.540 2.74 0.770 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.590 1.94 0.780 ;
        RECT 1.90 0.320 1.98 0.670 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.320 1.74 0.820 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.81 0.380 0.89 0.880 ;
        RECT 0.62 0.800 0.89 0.880 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.375 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.375 0.06 ;
    END
  END VSS
END MX3X2

MACRO MXI2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X2 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 0.260 1.91 0.400 ;
        RECT 1.86 0.340 1.92 0.980 ;
        RECT 1.86 0.400 1.94 0.530 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.500 1.54 0.910 ;
        RECT 1.46 0.500 1.62 0.720 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.69 0.500 0.77 0.750 ;
        RECT 0.44 0.590 0.77 0.750 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.750 0.34 0.910 ;
        RECT 0.86 0.640 0.93 0.910 ;
        RECT 0.28 0.850 0.93 0.910 ;
        RECT 1.14 0.500 1.20 0.700 ;
        RECT 0.86 0.640 1.20 0.700 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.835 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.835 0.06 ;
    END
  END VSS
END MXI2X2

MACRO MXI2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X6 0 0 ;
  SIZE 3.240 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.03 0.200 2.09 0.560 ;
        RECT 2.03 0.660 2.09 0.980 ;
        RECT 2.03 0.500 2.32 0.560 ;
        RECT 2.26 0.500 2.32 0.720 ;
        RECT 2.26 0.590 2.34 0.720 ;
        RECT 2.03 0.660 2.34 0.720 ;
        RECT 2.44 0.200 2.50 0.980 ;
        RECT 2.26 0.590 2.91 0.650 ;
        RECT 2.81 0.430 2.87 0.650 ;
        RECT 2.85 0.200 2.91 0.490 ;
        RECT 2.85 0.590 2.91 0.980 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.360 1.34 1.060 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.290 0.54 0.600 ;
        RECT 0.59 0.230 0.67 0.420 ;
        RECT 0.46 0.290 0.67 0.420 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.580 0.34 0.710 ;
        RECT 0.30 0.650 0.36 0.860 ;
        RECT 0.77 0.560 0.83 0.860 ;
        RECT 0.30 0.800 0.83 0.860 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.240 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.240 0.06 ;
    END
  END VSS
END MXI2X6

MACRO MXI4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X2 0 0 ;
  SIZE 5.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.31 0.260 4.72 0.350 ;
        RECT 4.64 0.260 4.72 0.720 ;
        RECT 4.64 0.490 4.74 0.620 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 0.400 1.92 0.950 ;
    END
  END C
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.250 0.34 0.520 ;
        RECT 0.26 0.250 0.73 0.330 ;
        RECT 0.65 0.250 0.73 0.460 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.15 0.400 1.26 0.950 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.530 0.54 0.940 ;
        RECT 0.46 0.760 0.73 0.840 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.31 0.480 3.37 0.910 ;
        RECT 3.39 0.390 3.45 0.540 ;
        RECT 3.31 0.480 3.45 0.540 ;
        RECT 4.96 0.430 5.02 0.910 ;
        RECT 3.31 0.850 5.02 0.910 ;
        RECT 5.04 0.370 5.17 0.500 ;
        RECT 4.96 0.430 5.17 0.500 ;
    END
  END S1
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.420 2.94 0.920 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.400 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.400 0.06 ;
    END
  END VSS
END MXI4X2


MACRO DFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX2 0 0 ;
  SIZE 4.995 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.300 3.74 0.530 ;
        RECT 3.66 0.350 3.90 0.400 ;
        RECT 3.84 0.230 3.90 0.980 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.330 3.34 0.980 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.330 2.94 0.830 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.640 0.36 0.970 ;
        RECT 0.23 0.900 0.36 0.970 ;
        RECT 0.37 0.400 0.45 0.710 ;
        RECT 0.28 0.640 0.45 0.710 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.995 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.995 0.06 ;
    END
  END VSS
END DFFX2

MACRO BUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX4 0 0 ;
  SIZE 1.620 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.220 0.29 0.840 ;
        RECT 0.28 0.160 0.34 0.280 ;
        RECT 0.26 0.780 0.34 0.980 ;
        RECT 0.26 0.780 0.34 0.910 ;
        RECT 0.23 0.780 0.76 0.840 ;
        RECT 0.23 0.220 0.72 0.280 ;
        RECT 0.70 0.780 0.76 0.980 ;
        RECT 0.67 0.200 0.79 0.260 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.96 0.580 1.04 0.950 ;
        RECT 1.05 0.440 1.13 0.660 ;
        RECT 0.96 0.580 1.13 0.660 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.620 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.620 0.06 ;
    END
  END VSS
END BUFX4

MACRO BUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX6 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.370 1.54 0.870 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 0.200 0.23 0.970 ;
        RECT 0.16 0.590 0.24 0.770 ;
        RECT 0.58 0.200 0.64 0.460 ;
        RECT 0.58 0.720 0.64 0.970 ;
        RECT 0.16 0.720 1.05 0.770 ;
        RECT 0.99 0.200 1.05 0.460 ;
        RECT 0.16 0.390 1.05 0.460 ;
        RECT 0.99 0.720 1.05 0.970 ;
    END
  END Y
END BUFX6

MACRO NAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X2 0 0 ;
  SIZE 1.215 BY 1.2 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.87 0.260 0.95 0.980 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.52 0.420 0.58 0.720 ;
        RECT 0.26 0.420 0.58 0.520 ;
        RECT 0.26 0.220 0.32 0.520 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.10 0.400 0.17 0.980 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.215 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.215 0.06 ;
    END
  END VSS
END NAND2X2

MACRO XOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X2 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.400 0.34 0.530 ;
        RECT 0.28 0.290 0.34 1.020 ;
        RECT 0.28 0.960 0.43 1.020 ;
        RECT 0.38 0.230 0.43 0.360 ;
        RECT 0.28 0.290 0.43 0.360 ;
        RECT 0.38 0.960 0.43 1.070 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.620 1.56 0.690 ;
        RECT 1.44 0.610 1.56 0.700 ;
        RECT 1.33 0.610 1.79 0.680 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.60 0.610 0.80 0.700 ;
        RECT 0.72 0.610 0.80 1.000 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS

END XOR2X2

MACRO XNOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X2 0 0 ;
  SIZE 2.565 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.340 0.54 0.920 ;
        RECT 0.42 0.840 0.54 0.920 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.59 0.610 2.09 0.700 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.490 0.91 0.700 ;
        RECT 0.64 0.610 1.01 0.700 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.565 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.565 0.06 ;
    END
  END VSS
END XNOR2X2

MACRO SDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX2 0 0 ;
  SIZE 5.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.590 0.36 0.720 ;
        RECT 0.30 0.340 0.36 0.980 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.20 0.300 4.25 0.680 ;
        RECT 4.44 0.300 4.56 0.470 ;
        RECT 5.03 0.610 5.17 0.680 ;
        RECT 4.20 0.300 5.14 0.360 ;
        RECT 5.08 0.300 5.14 0.700 ;
        RECT 5.04 0.610 5.17 0.700 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.84 0.460 4.92 0.770 ;
        RECT 4.66 0.590 4.92 0.770 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.300 3.74 0.530 ;
        RECT 3.66 0.450 3.94 0.530 ;
        RECT 3.85 0.450 3.94 0.810 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.740 0.54 0.910 ;
        RECT 0.74 0.490 0.81 0.820 ;
        RECT 0.46 0.740 0.81 0.820 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.400 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.400 0.06 ;
    END
  END VSS

END SDFFHQX2

MACRO SDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX8 0 0 ;
  SIZE 6.750 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.54 0.490 5.59 0.760 ;
        RECT 5.54 0.490 5.69 0.560 ;
        RECT 5.62 0.450 6.40 0.500 ;
        RECT 6.24 0.420 6.40 0.500 ;
        RECT 6.34 0.420 6.40 0.540 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.87 0.610 6.17 0.810 ;
        RECT 5.87 0.610 6.24 0.690 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.450 5.14 0.720 ;
        RECT 5.06 0.590 5.28 0.720 ;
        RECT 5.20 0.590 5.28 0.810 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.72 0.390 2.83 0.700 ;
        RECT 2.56 0.610 2.83 0.700 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.340 0.23 0.980 ;
        RECT 0.17 0.340 0.24 0.530 ;
        RECT 0.16 0.400 0.24 0.530 ;
        RECT 0.58 0.340 0.64 0.980 ;
        RECT 0.16 0.470 1.05 0.530 ;
        RECT 0.99 0.340 1.05 0.980 ;
        RECT 0.99 0.540 1.41 0.600 ;
        RECT 1.35 0.390 1.41 0.760 ;
        RECT 1.40 0.330 1.46 0.450 ;
        RECT 1.40 0.700 1.46 0.980 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 6.750 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 6.750 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal2 ;
        RECT 0.81 0.225 0.91 0.975 ;
        RECT 3.20 0.225 3.32 0.775 ;
        RECT 4.61 0.225 4.81 0.975 ;
        RECT 1.82 0.325 2.12 0.875 ;
  END
END SDFFHQX8

MACRO SDFFQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX2 0 0 ;
  SIZE 4.995 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.400 0.36 0.530 ;
        RECT 0.30 0.200 0.36 0.980 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.75 0.590 3.81 0.760 ;
        RECT 3.77 0.450 3.83 0.640 ;
        RECT 4.04 0.420 4.17 0.500 ;
        RECT 3.77 0.450 4.48 0.500 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.20 0.610 4.61 0.700 ;
        RECT 4.43 0.610 4.61 0.770 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.420 3.34 0.770 ;
        RECT 3.26 0.590 3.49 0.720 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.410 0.74 0.910 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.995 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.995 0.06 ;
    END
  END VSS
END SDFFQX2

MACRO SDFFQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX4 0 0 ;
  SIZE 5.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.51 0.450 4.58 0.780 ;
        RECT 4.46 0.730 4.58 0.780 ;
        RECT 5.04 0.420 5.17 0.500 ;
        RECT 4.51 0.450 5.17 0.500 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.83 0.610 4.94 0.810 ;
        RECT 4.83 0.610 5.21 0.700 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.00 0.560 4.17 0.700 ;
        RECT 4.08 0.560 4.17 0.780 ;
        RECT 4.00 0.560 4.36 0.680 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.450 0.31 0.770 ;
        RECT 0.26 0.300 0.34 0.530 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.400 0.57 0.530 ;
        RECT 0.51 0.370 0.57 0.980 ;
        RECT 0.48 0.370 0.60 0.460 ;
        RECT 0.46 0.400 0.94 0.460 ;
        RECT 0.88 0.370 0.94 0.740 ;
        RECT 0.92 0.690 0.98 0.980 ;
        RECT 0.88 0.370 1.07 0.430 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.400 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.400 0.06 ;
    END
  END VSS
END SDFFQX4

MACRO SDFFRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX8 0 0 ;
  SIZE 7.965 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.78 0.450 6.84 0.720 ;
        RECT 6.78 0.450 7.56 0.500 ;
        RECT 7.34 0.420 7.56 0.510 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.13 0.610 7.37 0.720 ;
        RECT 7.13 0.610 7.61 0.700 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.400 6.34 0.530 ;
        RECT 6.26 0.420 6.52 0.500 ;
        RECT 6.44 0.420 6.52 0.700 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.54 0.390 3.66 0.720 ;
        RECT 3.40 0.610 3.66 0.720 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.83 0.520 1.96 0.670 ;
        RECT 1.91 0.240 1.96 0.670 ;
        RECT 1.81 0.600 1.96 0.670 ;
        RECT 1.91 0.240 2.45 0.310 ;
        RECT 2.39 0.240 2.45 0.660 ;
        RECT 2.39 0.590 2.54 0.660 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.20 0.470 0.26 0.980 ;
        RECT 0.26 0.340 0.34 0.530 ;
        RECT 0.60 0.470 0.67 0.980 ;
        RECT 0.69 0.340 0.75 0.530 ;
        RECT 1.01 0.470 1.07 0.980 ;
        RECT 1.10 0.340 1.16 0.530 ;
        RECT 0.20 0.470 1.48 0.530 ;
        RECT 1.43 0.400 1.48 0.980 ;
        RECT 1.51 0.340 1.57 0.460 ;
        RECT 1.43 0.400 1.57 0.460 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 7.965 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 7.965 0.06 ;
    END
  END VSS
END SDFFRHQX8

MACRO SDFFRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX2 0 0 ;
  SIZE 6.615 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 0.290 1.14 0.790 ;
        RECT 1.05 0.400 1.14 0.530 ;
        RECT 1.05 0.710 1.18 0.790 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.290 0.73 0.790 ;
        RECT 0.56 0.710 0.73 0.790 ;
        RECT 0.65 0.400 0.74 0.530 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.63 0.400 5.71 0.680 ;
        RECT 5.63 0.400 6.14 0.480 ;
        RECT 6.06 0.400 6.14 0.530 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.81 0.580 5.89 0.880 ;
        RECT 5.63 0.800 5.89 0.880 ;
        RECT 5.81 0.580 5.94 0.660 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.590 5.14 0.820 ;
        RECT 5.13 0.400 5.21 0.670 ;
    END
  END SI
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.38 0.340 2.52 0.400 ;
        RECT 2.46 0.340 2.52 0.610 ;
        RECT 2.46 0.480 2.54 0.610 ;
        RECT 2.46 0.550 2.84 0.610 ;
        RECT 2.78 0.550 2.84 0.940 ;
        RECT 2.78 0.880 3.77 0.940 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.370 1.52 0.740 ;
        RECT 1.44 0.370 1.64 0.500 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 6.615 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 6.615 0.06 ;
    END
  END VSS
END SDFFRX2

MACRO SDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX2 0 0 ;
  SIZE 5.805 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.86 0.300 4.96 0.430 ;
        RECT 4.90 0.270 4.96 0.980 ;
        RECT 4.87 0.270 4.99 0.330 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.40 0.270 4.52 0.330 ;
        RECT 4.46 0.270 4.52 0.980 ;
        RECT 4.46 0.300 4.54 0.430 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.260 4.14 0.760 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.18 0.540 1.26 0.980 ;
        RECT 1.26 0.490 1.34 0.620 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.590 0.74 0.670 ;
        RECT 0.66 0.590 0.74 0.900 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.210 0.34 0.340 ;
        RECT 0.23 0.210 0.74 0.300 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.805 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.805 0.06 ;
    END
  END VSS
END SDFFX2

MACRO SDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX4 0 0 ;
  SIZE 5.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.47 0.610 4.53 0.730 ;
        RECT 4.50 0.460 4.56 0.670 ;
        RECT 5.04 0.420 5.17 0.510 ;
        RECT 4.50 0.460 5.17 0.510 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.82 0.610 5.06 0.780 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.590 3.94 0.720 ;
        RECT 3.86 0.640 4.21 0.720 ;
        RECT 4.13 0.550 4.21 0.730 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.490 0.34 0.990 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.590 0.54 0.870 ;
        RECT 0.53 0.340 0.58 0.650 ;
        RECT 1.00 0.340 1.06 0.870 ;
        RECT 0.46 0.810 1.06 0.870 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.400 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.400 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal2 ;
        RECT 3.00 0.225 3.32 0.775 ;
        RECT 1.22 0.225 1.72 0.975 ;
  END
END SDFFHQX4

MACRO OR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X2 0 0 ;
  SIZE 1.350 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.77 0.190 0.82 0.310 ;
        RECT 0.77 0.710 0.82 0.980 ;
        RECT 0.77 0.250 0.92 0.310 ;
        RECT 0.86 0.250 0.92 0.760 ;
        RECT 0.77 0.710 0.92 0.760 ;
        RECT 0.86 0.400 0.94 0.530 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 0.570 0.49 0.960 ;
        RECT 0.41 0.610 0.52 0.960 ;
        RECT 0.41 0.610 0.60 0.700 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.10 0.210 0.18 0.340 ;
        RECT 0.11 0.260 0.19 0.700 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.350 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.350 0.06 ;
    END
  END VSS
END OR2X2

MACRO NOR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X8 0 0 ;
  SIZE 3.375 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.790 0.71 0.990 ;
        RECT 1.30 0.790 1.36 0.990 ;
        RECT 2.19 0.790 2.25 0.990 ;
        RECT 0.66 0.790 3.14 0.850 ;
        RECT 2.92 0.760 2.98 0.990 ;
        RECT 0.32 0.290 3.14 0.350 ;
        RECT 3.08 0.290 3.14 0.910 ;
        RECT 2.92 0.760 3.14 0.910 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.69 0.610 0.91 0.670 ;
        RECT 1.41 0.610 1.53 0.700 ;
        RECT 2.02 0.610 2.15 0.700 ;
        RECT 2.63 0.610 2.93 0.660 ;
        RECT 0.85 0.630 2.77 0.700 ;
        RECT 2.71 0.600 2.93 0.660 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.580 0.54 0.640 ;
        RECT 0.48 0.450 0.54 0.720 ;
        RECT 0.46 0.580 0.54 0.720 ;
        RECT 1.01 0.450 1.13 0.530 ;
        RECT 1.81 0.450 1.93 0.530 ;
        RECT 0.48 0.450 2.31 0.510 ;
        RECT 2.25 0.480 2.56 0.530 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.375 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.375 0.06 ;
    END
  END VSS
END NOR2X8

MACRO OR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X4 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.97 0.650 1.03 0.980 ;
        RECT 0.94 0.200 1.06 0.260 ;
        RECT 1.01 0.220 1.52 0.280 ;
        RECT 0.97 0.650 1.52 0.720 ;
        RECT 1.40 0.160 1.46 0.280 ;
        RECT 1.40 0.810 1.46 0.980 ;
        RECT 1.46 0.220 1.52 0.870 ;
        RECT 1.46 0.400 1.54 0.530 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.60 0.540 0.74 0.660 ;
        RECT 0.66 0.540 0.74 0.990 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.10 0.400 0.18 0.630 ;
        RECT 0.10 0.400 0.34 0.480 ;
        RECT 0.27 0.400 0.34 0.740 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS
END OR2X4

MACRO NOR2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X6 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.230 0.34 0.360 ;
        RECT 0.58 0.820 0.64 0.980 ;
        RECT 0.69 0.230 0.74 0.360 ;
        RECT 1.09 0.230 1.16 0.360 ;
        RECT 1.23 0.820 1.28 0.980 ;
        RECT 1.50 0.230 1.56 0.360 ;
        RECT 1.92 0.230 1.98 0.360 ;
        RECT 1.92 0.820 1.98 0.980 ;
        RECT 0.28 0.290 2.38 0.360 ;
        RECT 2.26 0.780 2.34 0.910 ;
        RECT 2.32 0.290 2.38 0.880 ;
        RECT 0.58 0.820 2.38 0.880 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.61 0.610 0.83 0.680 ;
        RECT 1.16 0.610 1.27 0.720 ;
        RECT 0.78 0.650 1.89 0.720 ;
        RECT 1.83 0.610 2.06 0.700 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.21 0.590 0.34 0.650 ;
        RECT 0.28 0.460 0.34 0.720 ;
        RECT 0.26 0.590 0.34 0.720 ;
        RECT 0.94 0.460 1.05 0.560 ;
        RECT 1.55 0.460 1.67 0.560 ;
        RECT 0.28 0.460 2.22 0.510 ;
        RECT 2.16 0.460 2.22 0.680 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.835 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.835 0.06 ;
    END
  END VSS
END NOR2X6

MACRO NOR2BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX4 0 0 ;
  SIZE 2.430 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.10 0.290 0.16 0.850 ;
        RECT 0.10 0.610 0.22 0.700 ;
        RECT 0.28 0.230 0.34 0.350 ;
        RECT 0.54 0.790 0.59 0.980 ;
        RECT 0.69 0.230 0.74 0.350 ;
        RECT 0.10 0.790 1.22 0.850 ;
        RECT 1.09 0.230 1.16 0.350 ;
        RECT 1.16 0.790 1.22 0.980 ;
        RECT 1.50 0.230 1.56 0.350 ;
        RECT 0.10 0.290 1.56 0.350 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.610 1.25 0.700 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.780 1.54 0.910 ;
        RECT 1.69 0.610 1.77 0.860 ;
        RECT 1.46 0.780 1.77 0.860 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.430 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.430 0.06 ;
    END
  END VSS
END NOR2BX4

MACRO NOR3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X8 0 0 ;
  SIZE 5.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.00 0.890 1.06 0.980 ;
        RECT 2.25 0.890 2.31 0.980 ;
        RECT 3.77 0.890 3.83 0.980 ;
        RECT 1.00 0.890 4.97 0.950 ;
        RECT 4.91 0.700 4.97 0.980 ;
        RECT 5.03 0.200 5.08 0.880 ;
        RECT 4.91 0.700 5.08 0.880 ;
        RECT 4.91 0.800 5.17 0.880 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.31 0.530 0.37 0.700 ;
        RECT 0.23 0.610 0.37 0.700 ;
        RECT 0.23 0.630 0.57 0.700 ;
        RECT 0.52 0.630 0.57 0.790 ;
        RECT 1.62 0.570 1.75 0.630 ;
        RECT 1.69 0.570 1.75 0.790 ;
        RECT 2.83 0.570 2.89 0.790 ;
        RECT 2.83 0.570 2.95 0.630 ;
        RECT 4.19 0.570 4.25 0.790 ;
        RECT 0.52 0.730 4.25 0.790 ;
        RECT 4.19 0.570 4.31 0.630 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.480 0.73 0.530 ;
        RECT 0.68 0.480 0.73 0.630 ;
        RECT 1.21 0.420 1.27 0.630 ;
        RECT 0.68 0.570 1.27 0.630 ;
        RECT 1.21 0.420 1.32 0.480 ;
        RECT 1.91 0.410 1.97 0.530 ;
        RECT 1.27 0.410 2.19 0.470 ;
        RECT 2.12 0.410 2.19 0.630 ;
        RECT 2.56 0.420 2.62 0.630 ;
        RECT 2.12 0.570 2.62 0.630 ;
        RECT 2.56 0.420 2.68 0.480 ;
        RECT 2.62 0.410 3.29 0.470 ;
        RECT 3.23 0.420 3.59 0.480 ;
        RECT 3.54 0.420 3.59 0.630 ;
        RECT 3.92 0.420 3.98 0.630 ;
        RECT 3.54 0.570 3.98 0.630 ;
        RECT 3.92 0.420 4.09 0.480 ;
        RECT 4.03 0.410 4.47 0.470 ;
        RECT 4.41 0.420 4.76 0.490 ;
        RECT 4.63 0.420 4.76 0.500 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.83 0.230 1.07 0.470 ;
        RECT 2.34 0.230 2.41 0.470 ;
        RECT 2.29 0.410 2.41 0.470 ;
        RECT 3.69 0.230 3.75 0.470 ;
        RECT 3.69 0.410 3.81 0.470 ;
        RECT 0.83 0.230 4.92 0.290 ;
        RECT 4.87 0.230 4.92 0.520 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.400 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.400 0.06 ;
    END
  END VSS
END NOR3X8

MACRO NAND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X6 0 0 ;
  SIZE 2.97 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 0.810 0.47 0.980 ;
        RECT 0.64 0.230 0.70 0.360 ;
        RECT 0.81 0.810 0.88 0.980 ;
        RECT 1.23 0.810 1.29 0.980 ;
        RECT 1.54 0.230 1.60 0.360 ;
        RECT 1.65 0.810 1.71 0.980 ;
        RECT 2.06 0.810 2.12 0.980 ;
        RECT 2.16 0.230 2.22 0.360 ;
        RECT 0.41 0.810 2.76 0.870 ;
        RECT 2.46 0.810 2.52 0.980 ;
        RECT 0.64 0.290 2.76 0.360 ;
        RECT 2.66 0.780 2.74 0.910 ;
        RECT 2.70 0.290 2.76 0.880 ;
        RECT 2.46 0.810 2.76 0.880 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.71 0.610 0.97 0.680 ;
        RECT 1.45 0.610 1.56 0.720 ;
        RECT 0.92 0.650 2.08 0.720 ;
        RECT 2.04 0.610 2.19 0.700 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.400 0.54 0.560 ;
        RECT 0.34 0.490 0.54 0.560 ;
        RECT 1.07 0.460 1.20 0.560 ;
        RECT 1.75 0.460 1.88 0.540 ;
        RECT 0.46 0.460 2.60 0.510 ;
        RECT 2.54 0.460 2.60 0.680 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.97 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.97 0.06 ;
    END
  END VSS

END NAND2X6


MACRO NAND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X4 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 0.790 0.40 0.980 ;
        RECT 0.63 0.270 0.75 0.340 ;
        RECT 0.75 0.790 0.81 0.980 ;
        RECT 1.16 0.790 1.22 0.980 ;
        RECT 1.25 0.270 1.37 0.360 ;
        RECT 1.57 0.790 1.63 0.980 ;
        RECT 0.70 0.290 1.77 0.360 ;
        RECT 1.64 0.610 1.77 0.700 ;
        RECT 1.71 0.290 1.77 0.850 ;
        RECT 0.34 0.790 1.77 0.850 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.610 1.29 0.700 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.420 0.36 0.510 ;
        RECT 0.23 0.460 1.60 0.510 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS
END NAND2X4

MACRO NAND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X8 0 0 ;
  SIZE 3.375 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.690 0.35 0.980 ;
        RECT 0.70 0.750 0.77 0.980 ;
        RECT 1.11 0.750 1.18 0.980 ;
        RECT 1.52 0.750 1.58 0.980 ;
        RECT 1.94 0.750 2.00 0.980 ;
        RECT 2.34 0.750 2.41 0.980 ;
        RECT 2.75 0.750 2.81 0.980 ;
        RECT 0.47 0.250 3.14 0.300 ;
        RECT 3.06 0.680 3.14 0.810 ;
        RECT 3.08 0.250 3.14 0.810 ;
        RECT 0.29 0.750 3.14 0.810 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.54 0.560 0.81 0.630 ;
        RECT 1.43 0.560 1.55 0.650 ;
        RECT 2.04 0.560 2.17 0.650 ;
        RECT 2.63 0.510 2.77 0.650 ;
        RECT 0.75 0.590 2.77 0.650 ;
        RECT 2.63 0.510 2.88 0.580 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.320 0.36 0.490 ;
        RECT 0.91 0.400 1.03 0.490 ;
        RECT 1.77 0.400 1.90 0.490 ;
        RECT 0.23 0.400 2.33 0.470 ;
        RECT 2.27 0.430 2.51 0.490 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.375 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.375 0.06 ;
    END
  END VSS
END NAND2X8

MACRO NOR4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X2 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.250 0.40 0.310 ;
        RECT 0.71 0.250 0.83 0.330 ;
        RECT 1.16 0.250 1.27 0.330 ;
        RECT 1.59 0.250 1.71 0.330 ;
        RECT 0.34 0.270 1.94 0.330 ;
        RECT 1.88 0.270 1.94 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.620 0.32 0.990 ;
        RECT 1.66 0.780 1.74 0.990 ;
        RECT 1.68 0.620 1.74 0.990 ;
        RECT 0.26 0.920 1.74 0.990 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 0.630 0.54 0.700 ;
        RECT 0.46 0.590 0.54 0.720 ;
        RECT 0.48 0.590 0.54 0.820 ;
        RECT 1.44 0.640 1.50 0.820 ;
        RECT 0.48 0.760 1.50 0.820 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.27 0.420 1.33 0.660 ;
        RECT 0.64 0.610 1.33 0.660 ;
        RECT 1.27 0.420 1.56 0.500 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.420 1.14 0.500 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS
END NOR4X2


MACRO NAND3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X8 0 0 ;
  SIZE 4.995 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.71 0.860 3.77 0.980 ;
        RECT 3.71 0.910 4.17 0.980 ;
        RECT 4.12 0.810 4.17 0.980 ;
        RECT 4.46 0.780 4.62 0.910 ;
        RECT 4.12 0.850 4.62 0.910 ;
        RECT 0.48 0.210 4.62 0.270 ;
        RECT 4.56 0.210 4.62 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.590 0.34 0.720 ;
        RECT 0.28 0.590 0.34 0.890 ;
        RECT 0.28 0.830 0.54 0.890 ;
        RECT 1.28 0.690 1.34 0.910 ;
        RECT 0.47 0.850 1.34 0.910 ;
        RECT 1.28 0.690 1.40 0.760 ;
        RECT 1.28 0.700 1.80 0.760 ;
        RECT 1.74 0.700 1.80 0.910 ;
        RECT 2.55 0.690 2.67 0.740 ;
        RECT 2.61 0.690 2.67 0.910 ;
        RECT 3.54 0.700 3.60 0.910 ;
        RECT 1.74 0.850 3.60 0.910 ;
        RECT 3.54 0.700 3.79 0.760 ;
        RECT 3.73 0.690 3.86 0.740 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 0.680 0.69 0.740 ;
        RECT 1.04 0.520 1.10 0.750 ;
        RECT 0.64 0.690 1.10 0.750 ;
        RECT 1.04 0.520 1.56 0.590 ;
        RECT 1.50 0.540 1.96 0.600 ;
        RECT 1.90 0.540 1.96 0.750 ;
        RECT 2.28 0.540 2.34 0.750 ;
        RECT 1.90 0.690 2.34 0.750 ;
        RECT 2.28 0.540 2.40 0.600 ;
        RECT 2.34 0.520 2.83 0.590 ;
        RECT 2.77 0.540 3.03 0.600 ;
        RECT 2.97 0.540 3.03 0.750 ;
        RECT 3.38 0.540 3.44 0.750 ;
        RECT 2.97 0.690 3.44 0.750 ;
        RECT 3.38 0.540 3.63 0.600 ;
        RECT 3.51 0.520 4.25 0.590 ;
        RECT 4.04 0.520 4.25 0.700 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.400 0.94 0.590 ;
        RECT 0.80 0.530 0.94 0.590 ;
        RECT 2.06 0.360 2.12 0.590 ;
        RECT 2.06 0.530 2.18 0.590 ;
        RECT 3.23 0.360 3.29 0.590 ;
        RECT 3.17 0.530 3.29 0.590 ;
        RECT 0.88 0.360 4.41 0.420 ;
        RECT 4.34 0.360 4.41 0.600 ;
        RECT 4.34 0.540 4.46 0.600 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.995 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.995 0.06 ;
    END
  END VSS

END NAND3X8

MACRO NOR3BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX2 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.200 0.14 0.720 ;
        RECT 0.06 0.590 0.14 0.720 ;
        RECT 0.06 0.660 0.90 0.720 ;
        RECT 0.83 0.660 0.90 0.980 ;
        RECT 0.08 0.200 1.50 0.260 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 0.600 1.14 0.680 ;
        RECT 1.06 0.600 1.14 0.980 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 0.440 1.34 0.500 ;
        RECT 1.26 0.440 1.34 0.720 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.60 0.440 1.68 0.880 ;
        RECT 1.60 0.440 1.74 0.720 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS
END NOR3BX2

MACRO OA21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X2 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.20 0.470 1.26 0.980 ;
        RECT 1.26 0.400 1.34 0.530 ;
        RECT 1.28 0.370 1.50 0.430 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.360 0.34 0.860 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.590 0.54 0.730 ;
        RECT 0.62 0.390 0.70 0.660 ;
        RECT 0.46 0.590 0.70 0.660 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.200 0.94 0.620 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS
END OA21X2

MACRO OAI221X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X2 0 0 ;
  SIZE 2.97 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.44 0.270 2.50 0.980 ;
        RECT 0.66 0.920 2.50 0.980 ;
        RECT 2.44 0.590 2.54 0.720 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.490 0.34 0.620 ;
        RECT 0.22 0.560 0.34 0.620 ;
        RECT 0.28 0.490 0.34 0.750 ;
        RECT 0.94 0.540 1.00 0.750 ;
        RECT 0.28 0.690 1.00 0.750 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.40 0.540 1.46 0.750 ;
        RECT 2.06 0.490 2.14 0.750 ;
        RECT 1.40 0.690 2.14 0.750 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.410 0.71 0.500 ;
        RECT 0.64 0.410 0.71 0.600 ;
        RECT 0.64 0.510 0.84 0.600 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.69 0.410 1.77 0.600 ;
        RECT 1.56 0.510 1.77 0.600 ;
        RECT 1.69 0.410 1.96 0.500 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.260 2.34 0.750 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.97 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.97 0.06 ;
    END
  END VSS

END OAI221X2

MACRO OAI222X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X2 0 0 ;
  SIZE 3.645 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.42 0.210 2.48 0.360 ;
        RECT 2.83 0.210 2.88 0.360 ;
        RECT 2.42 0.290 3.32 0.360 ;
        RECT 3.26 0.290 3.32 0.980 ;
        RECT 0.62 0.920 3.32 0.980 ;
        RECT 3.26 0.400 3.34 0.530 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.640 0.34 0.850 ;
        RECT 0.86 0.590 0.94 0.850 ;
        RECT 0.28 0.790 0.94 0.850 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.42 0.630 1.54 0.700 ;
        RECT 1.46 0.590 1.54 0.850 ;
        RECT 2.08 0.640 2.14 0.850 ;
        RECT 1.46 0.790 2.14 0.850 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.640 2.32 0.850 ;
        RECT 2.86 0.590 2.92 0.850 ;
        RECT 2.26 0.790 2.92 0.850 ;
        RECT 2.86 0.590 2.94 0.720 ;
        RECT 2.86 0.590 2.98 0.650 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.480 0.65 0.700 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 0.460 2.76 0.700 ;
        RECT 2.42 0.580 2.76 0.700 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 0.460 1.98 0.530 ;
        RECT 1.83 0.460 1.98 0.700 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.645 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.645 0.06 ;
    END
  END VSS

END OAI222X2

MACRO OAI2BB1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X4 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.12 0.390 0.17 0.980 ;
        RECT 0.06 0.780 0.17 0.980 ;
        RECT 0.51 0.370 0.63 0.450 ;
        RECT 0.12 0.390 1.15 0.450 ;
        RECT 1.09 0.370 1.36 0.430 ;
        RECT 0.06 0.920 1.64 0.980 ;
    END
  END Y
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.79 0.420 1.96 0.500 ;
        RECT 1.89 0.420 1.96 0.700 ;
        RECT 1.89 0.620 2.10 0.700 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.36 0.560 2.44 0.860 ;
        RECT 2.36 0.780 2.54 0.860 ;
        RECT 2.46 0.780 2.54 0.960 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.550 0.54 0.720 ;
        RECT 0.28 0.550 1.69 0.610 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.835 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.835 0.06 ;
    END
  END VSS

END OAI2BB1X4

MACRO OAI31X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X2 0 0 ;
  SIZE 2.430 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.680 1.54 0.980 ;
        RECT 1.46 0.750 1.71 0.980 ;
        RECT 0.91 0.890 1.71 0.980 ;
        RECT 1.66 0.750 1.71 0.980 ;
        RECT 1.70 0.250 1.76 0.810 ;
        RECT 1.70 0.250 1.88 0.300 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 0.620 1.17 0.780 ;
        RECT 0.89 0.700 1.17 0.780 ;
        RECT 0.94 0.620 1.30 0.690 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.460 0.74 0.620 ;
        RECT 0.49 0.460 1.23 0.510 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 0.290 0.40 0.500 ;
        RECT 0.34 0.290 1.46 0.360 ;
        RECT 1.40 0.300 1.54 0.520 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.400 1.94 0.980 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.430 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.430 0.06 ;
    END
  END VSS
END OAI31X2

MACRO OR4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X6 0 0 ;
  SIZE 3.375 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.00 0.780 2.06 0.980 ;
        RECT 2.09 0.200 2.15 0.380 ;
        RECT 2.00 0.780 2.74 0.840 ;
        RECT 2.41 0.780 2.47 0.980 ;
        RECT 2.50 0.200 2.56 0.380 ;
        RECT 2.66 0.330 2.72 0.910 ;
        RECT 2.41 0.780 2.74 0.910 ;
        RECT 2.41 0.850 2.88 0.910 ;
        RECT 2.82 0.850 2.88 0.980 ;
        RECT 2.91 0.200 2.97 0.380 ;
        RECT 2.09 0.330 2.97 0.380 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.30 0.490 0.36 0.980 ;
        RECT 1.66 0.410 1.72 0.980 ;
        RECT 0.30 0.900 1.72 0.980 ;
        RECT 1.66 0.580 1.74 0.710 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.390 0.54 0.670 ;
        RECT 0.46 0.520 0.58 0.670 ;
        RECT 1.50 0.490 1.56 0.670 ;
        RECT 0.46 0.610 1.56 0.670 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.220 1.36 0.300 ;
        RECT 1.30 0.220 1.36 0.510 ;
        RECT 0.68 0.450 1.36 0.510 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 0.220 0.96 0.350 ;
        RECT 0.68 0.270 1.14 0.350 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.375 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.375 0.06 ;
    END
  END VSS
END OR4X6

#### OLD MACROS

MACRO OA22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X2 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.470 1.50 0.980 ;
        RECT 1.46 0.370 1.54 0.530 ;
        RECT 1.46 0.370 1.61 0.430 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.00 0.780 1.08 0.970 ;
        RECT 1.00 0.780 1.34 0.860 ;
        RECT 1.26 0.780 1.34 0.910 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.480 0.54 0.980 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.480 0.34 0.980 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.480 0.74 0.980 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS

END OA22X2




MACRO TLATNTSCAX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX16 0 0 ;
  SIZE 7.830 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.62 0.300 4.67 0.420 ;
        RECT 4.66 0.360 4.72 0.980 ;
        RECT 4.66 0.590 4.74 0.720 ;
        RECT 5.00 0.370 5.12 0.430 ;
        RECT 5.07 0.610 5.13 0.980 ;
        RECT 5.07 0.380 5.50 0.450 ;
        RECT 5.43 0.330 5.50 0.680 ;
        RECT 5.48 0.610 5.54 0.980 ;
        RECT 5.81 0.370 5.94 0.430 ;
        RECT 5.89 0.610 5.95 0.980 ;
        RECT 5.89 0.380 6.32 0.450 ;
        RECT 6.25 0.330 6.32 0.680 ;
        RECT 6.30 0.610 6.36 0.980 ;
        RECT 6.63 0.370 6.75 0.430 ;
        RECT 6.71 0.610 6.77 0.980 ;
        RECT 6.71 0.380 7.13 0.450 ;
        RECT 4.66 0.610 7.18 0.680 ;
        RECT 7.08 0.330 7.13 0.680 ;
        RECT 7.12 0.610 7.18 0.980 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.250 0.74 0.750 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.250 0.54 0.750 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.340 0.14 0.750 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 7.830 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 7.830 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal2 ;
        RECT 0.90 0.225 1.00 0.975 ;
        RECT 3.20 0.225 3.32 0.775 ;
        RECT 4.71 0.225 4.81 0.975 ;
        RECT 6.71 0.325 6.81 0.875 ;
        RECT 1.82 0.325 1.92 0.875 ;
  END

END TLATNTSCAX16




MACRO AOI221X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X2 0 0 ;
  SIZE 2.97 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.590 1.14 0.720 ;
        RECT 1.08 0.250 1.14 0.850 ;
        RECT 0.60 0.250 2.17 0.310 ;
        RECT 1.08 0.790 2.28 0.850 ;
        RECT 2.22 0.790 2.28 0.940 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.610 1.94 0.700 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.580 0.74 0.880 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.420 0.36 0.510 ;
        RECT 0.28 0.410 0.96 0.490 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 0.420 1.77 0.510 ;
        RECT 1.24 0.440 1.94 0.510 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.06 0.610 2.56 0.700 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.97 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.97 0.06 ;
    END
  END VSS

END AOI221X2



MACRO NAND3BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX2 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.15 0.140 0.21 0.880 ;
        RECT 0.15 0.800 0.43 0.880 ;
        RECT 0.37 0.800 0.43 0.980 ;
        RECT 0.15 0.140 0.82 0.200 ;
        RECT 0.79 0.860 0.85 0.980 ;
        RECT 0.37 0.860 1.26 0.920 ;
        RECT 1.20 0.820 1.26 0.980 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.53 0.610 0.96 0.700 ;
        RECT 0.88 0.610 0.96 0.760 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.460 1.13 0.510 ;
        RECT 1.06 0.510 1.14 0.720 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.590 1.54 0.920 ;
        RECT 1.49 0.460 1.57 0.720 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS

END NAND3BX2


MACRO OR3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X2 0 0 ;
  SIZE 1.62 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.93 0.710 0.99 0.980 ;
        RECT 1.02 0.170 1.08 0.770 ;
        RECT 0.93 0.710 1.08 0.770 ;
        RECT 1.26 0.400 1.34 0.530 ;
        RECT 1.02 0.470 1.34 0.530 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.62 0.420 0.74 0.860 ;
        RECT 0.62 0.420 0.77 0.500 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.440 0.34 0.720 ;
        RECT 0.28 0.590 0.36 0.910 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.410 0.14 0.910 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.62 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.62 0.06 ;
    END
  END VSS

END OR3X2






MACRO AOI2BB2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X2 0 0 ;
  SIZE 3.240 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.41 0.250 1.67 0.310 ;
        RECT 1.86 0.590 1.94 0.720 ;
        RECT 1.88 0.270 1.94 0.850 ;
        RECT 2.10 0.790 2.16 0.940 ;
        RECT 1.61 0.270 2.33 0.330 ;
        RECT 2.27 0.250 2.40 0.310 ;
        RECT 1.88 0.790 2.57 0.850 ;
        RECT 2.51 0.790 2.57 0.940 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.08 0.610 2.56 0.700 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.04 0.420 2.63 0.500 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.400 0.54 0.900 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.260 0.34 0.760 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.240 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.240 0.06 ;
    END
  END VSS

END AOI2BB2X2

MACRO SEDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX2 0 0 ;
  SIZE 8.370 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.86 0.400 5.07 0.530 ;
        RECT 4.99 0.320 5.07 0.820 ;
        RECT 4.99 0.320 5.19 0.400 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.54 0.690 4.62 0.820 ;
        RECT 4.60 0.320 4.68 0.790 ;
        RECT 4.54 0.690 4.69 0.790 ;
        RECT 4.60 0.320 4.72 0.400 ;
        RECT 4.60 0.590 4.74 0.720 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.83 0.410 7.96 0.860 ;
        RECT 7.83 0.610 7.96 0.860 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.50 0.580 7.58 0.700 ;
        RECT 7.04 0.610 7.58 0.700 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.76 0.610 6.03 0.930 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.480 4.34 0.980 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.19 0.710 0.67 0.800 ;
        RECT 0.19 0.710 0.68 0.800 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.520 0.43 0.600 ;
        RECT 0.64 0.200 0.69 0.600 ;
        RECT 0.23 0.550 0.84 0.600 ;
        RECT 0.64 0.200 1.16 0.260 ;
        RECT 1.10 0.200 1.16 0.750 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 8.370 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 8.370 0.06 ;
    END
  END VSS

END SEDFFTRX2





MACRO OR4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X4 0 0 ;
  SIZE 2.430 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.39 0.790 1.45 0.980 ;
        RECT 1.44 0.210 1.50 0.350 ;
        RECT 1.39 0.790 1.94 0.850 ;
        RECT 1.79 0.790 1.85 0.980 ;
        RECT 1.85 0.210 1.94 0.350 ;
        RECT 1.44 0.280 1.94 0.350 ;
        RECT 1.88 0.210 1.94 0.980 ;
        RECT 1.79 0.790 1.94 0.980 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.590 0.74 0.940 ;
        RECT 0.67 0.450 0.74 0.720 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.450 0.56 0.920 ;
        RECT 0.46 0.600 0.56 0.920 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.410 0.34 0.910 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.280 1.34 0.530 ;
        RECT 1.00 0.450 1.34 0.530 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.430 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.430 0.06 ;
    END
  END VSS

END OR4X4


MACRO NAND3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X2 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.850 0.43 0.980 ;
        RECT 0.78 0.850 0.84 0.980 ;
        RECT 1.19 0.850 1.25 0.980 ;
        RECT 0.80 0.140 1.56 0.200 ;
        RECT 1.44 0.800 1.56 0.910 ;
        RECT 1.50 0.140 1.56 0.910 ;
        RECT 0.36 0.850 1.56 0.910 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.52 0.610 0.77 0.750 ;
        RECT 0.52 0.610 0.96 0.700 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.460 1.14 0.510 ;
        RECT 1.06 0.460 1.14 0.720 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.31 0.290 0.37 0.530 ;
        RECT 0.26 0.400 0.37 0.530 ;
        RECT 0.31 0.290 1.30 0.360 ;
        RECT 1.24 0.290 1.30 0.530 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS

END NAND3X2


MACRO NAND3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X4 0 0 ;
  SIZE 2.97 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 0.810 0.47 0.980 ;
        RECT 0.82 0.920 0.89 0.980 ;
        RECT 1.23 0.920 1.29 0.980 ;
        RECT 1.65 0.920 1.71 0.980 ;
        RECT 2.06 0.920 2.12 0.980 ;
        RECT 0.41 0.920 2.52 0.980 ;
        RECT 2.46 0.840 2.52 0.980 ;
        RECT 0.90 0.210 2.74 0.270 ;
        RECT 2.66 0.780 2.74 0.910 ;
        RECT 2.68 0.210 2.74 0.910 ;
        RECT 2.46 0.850 2.74 0.910 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.610 0.36 0.700 ;
        RECT 0.30 0.650 0.70 0.720 ;
        RECT 0.64 0.650 0.70 0.820 ;
        RECT 1.48 0.690 1.59 0.820 ;
        RECT 2.31 0.680 2.37 0.820 ;
        RECT 0.64 0.760 2.37 0.820 ;
        RECT 2.50 0.620 2.56 0.740 ;
        RECT 2.31 0.680 2.56 0.740 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.52 0.490 0.86 0.560 ;
        RECT 0.80 0.490 0.86 0.660 ;
        RECT 1.27 0.520 1.32 0.660 ;
        RECT 0.80 0.610 1.32 0.660 ;
        RECT 1.27 0.520 1.75 0.590 ;
        RECT 1.69 0.520 1.75 0.660 ;
        RECT 2.15 0.490 2.21 0.660 ;
        RECT 1.69 0.610 2.21 0.660 ;
        RECT 2.26 0.400 2.34 0.540 ;
        RECT 2.26 0.420 2.40 0.540 ;
        RECT 2.15 0.490 2.40 0.540 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.03 0.360 1.17 0.500 ;
        RECT 0.96 0.450 1.17 0.500 ;
        RECT 1.03 0.360 1.92 0.420 ;
        RECT 1.85 0.360 1.92 0.500 ;
        RECT 1.85 0.450 1.98 0.500 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.97 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.97 0.06 ;
    END
  END VSS

END NAND3X4



















MACRO ADDHX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX2 0 0 ;
  SIZE 3.240 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.21 0.330 2.34 0.400 ;
        RECT 2.26 0.330 2.34 0.790 ;
        RECT 2.26 0.710 2.41 0.790 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.77 0.360 1.14 0.440 ;
        RECT 1.06 0.360 1.14 0.850 ;
        RECT 0.86 0.790 1.14 0.850 ;
    END
  END CO
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.51 0.600 0.67 0.780 ;
        RECT 0.60 0.600 0.67 0.990 ;
        RECT 0.60 0.930 1.36 0.990 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.160 0.32 0.630 ;
        RECT 0.26 0.400 0.34 0.630 ;
        RECT 1.46 0.160 1.52 0.760 ;
        RECT 0.26 0.160 2.79 0.220 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.240 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.240 0.06 ;
    END
  END VSS

END ADDHX2








MACRO NOR2BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX2 0 0 ;
  SIZE 1.755 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.280 0.14 0.720 ;
        RECT 0.06 0.590 0.14 0.720 ;
        RECT 0.49 0.260 0.61 0.340 ;
        RECT 0.06 0.660 0.76 0.720 ;
        RECT 0.70 0.660 0.76 0.980 ;
        RECT 0.08 0.280 0.98 0.340 ;
        RECT 0.93 0.260 1.05 0.320 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.780 1.14 0.940 ;
        RECT 1.22 0.600 1.30 0.860 ;
        RECT 1.06 0.780 1.30 0.860 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.600 0.94 0.980 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.755 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.755 0.06 ;
    END
  END VSS

END NOR2BX2

MACRO AOI21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X4 0 0 ;
  SIZE 3.240 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.79 0.250 0.91 0.310 ;
        RECT 1.41 0.250 1.52 0.330 ;
        RECT 1.89 0.270 1.95 0.700 ;
        RECT 1.95 0.210 2.01 0.330 ;
        RECT 1.89 0.610 2.17 0.700 ;
        RECT 2.06 0.610 2.17 0.870 ;
        RECT 0.85 0.270 2.40 0.330 ;
        RECT 2.34 0.250 2.46 0.310 ;
        RECT 2.06 0.750 2.53 0.810 ;
        RECT 2.47 0.750 2.53 0.870 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.71 0.610 1.45 0.700 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.54 0.460 1.74 0.510 ;
        RECT 1.66 0.460 1.74 0.720 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.23 0.420 2.37 0.510 ;
        RECT 2.05 0.440 2.54 0.510 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.240 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.240 0.06 ;
    END
  END VSS

END AOI21X4

MACRO OR2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X6 0 0 ;
  SIZE 2.565 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.760 1.28 0.980 ;
        RECT 1.30 0.150 1.36 0.460 ;
        RECT 1.64 0.760 1.69 0.980 ;
        RECT 1.71 0.150 1.77 0.460 ;
        RECT 1.86 0.400 1.92 0.820 ;
        RECT 1.86 0.400 1.94 0.530 ;
        RECT 1.23 0.760 2.10 0.820 ;
        RECT 2.04 0.760 2.10 0.980 ;
        RECT 2.12 0.150 2.18 0.460 ;
        RECT 1.30 0.400 2.18 0.460 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.710 0.54 0.980 ;
        RECT 0.46 0.710 0.67 0.790 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.570 0.34 0.720 ;
        RECT 0.26 0.570 0.36 0.650 ;
        RECT 0.28 0.530 0.96 0.610 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.565 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.565 0.06 ;
    END
  END VSS

END OR2X6

MACRO OAI22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X2 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.820 0.70 0.980 ;
        RECT 0.94 0.420 0.99 0.880 ;
        RECT 0.83 0.800 0.99 0.880 ;
        RECT 1.10 0.250 1.16 0.490 ;
        RECT 0.94 0.420 1.16 0.490 ;
        RECT 1.10 0.250 1.25 0.360 ;
        RECT 0.64 0.820 1.47 0.880 ;
        RECT 1.41 0.820 1.47 0.980 ;
        RECT 1.10 0.290 1.58 0.360 ;
        RECT 1.52 0.250 1.66 0.310 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.610 0.34 0.910 ;
        RECT 0.26 0.610 0.66 0.690 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.630 1.74 0.720 ;
        RECT 1.66 0.630 1.74 0.910 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.20 0.420 0.83 0.500 ;
        RECT 0.76 0.420 0.83 0.540 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 0.590 1.34 0.660 ;
        RECT 1.26 0.460 1.34 0.720 ;
        RECT 1.26 0.460 1.73 0.530 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS

END OAI22X2




MACRO NOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X4 0 0 ;
  SIZE 2.430 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.230 0.49 0.360 ;
        RECT 0.74 0.790 0.80 0.980 ;
        RECT 0.84 0.230 0.91 0.360 ;
        RECT 1.25 0.230 1.31 0.360 ;
        RECT 1.41 0.790 1.47 0.980 ;
        RECT 1.67 0.230 1.73 0.360 ;
        RECT 0.43 0.290 1.96 0.360 ;
        RECT 1.83 0.610 1.96 0.700 ;
        RECT 1.91 0.290 1.96 0.850 ;
        RECT 0.74 0.790 1.96 0.850 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 0.610 1.42 0.700 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.460 0.54 0.720 ;
        RECT 0.36 0.460 1.79 0.510 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.430 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.430 0.06 ;
    END
  END VSS

END NOR2X4



MACRO NOR4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X8 0 0 ;
  SIZE 6.345 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.260 0.38 0.320 ;
        RECT 0.67 0.260 0.79 0.330 ;
        RECT 1.08 0.260 1.20 0.330 ;
        RECT 1.49 0.260 1.61 0.330 ;
        RECT 1.95 0.260 2.07 0.330 ;
        RECT 2.36 0.260 2.48 0.330 ;
        RECT 2.77 0.260 2.89 0.330 ;
        RECT 3.18 0.260 3.30 0.330 ;
        RECT 3.59 0.260 3.71 0.330 ;
        RECT 4.00 0.260 4.12 0.330 ;
        RECT 4.41 0.260 4.53 0.330 ;
        RECT 4.64 0.790 4.71 0.980 ;
        RECT 4.82 0.260 4.94 0.330 ;
        RECT 5.05 0.790 5.12 0.980 ;
        RECT 5.23 0.260 5.35 0.330 ;
        RECT 5.30 0.610 5.53 0.850 ;
        RECT 4.64 0.790 5.53 0.850 ;
        RECT 5.46 0.590 5.53 0.980 ;
        RECT 5.30 0.610 5.54 0.720 ;
        RECT 5.49 0.270 5.55 0.680 ;
        RECT 5.67 0.210 5.73 0.330 ;
        RECT 0.34 0.270 5.73 0.330 ;
        RECT 5.30 0.610 5.94 0.680 ;
        RECT 5.88 0.610 5.94 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.550 0.94 0.720 ;
        RECT 0.95 0.510 1.03 0.630 ;
        RECT 0.40 0.550 1.03 0.630 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.04 0.570 2.17 0.700 ;
        RECT 1.89 0.570 2.54 0.650 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.32 0.570 4.34 0.630 ;
        RECT 4.22 0.510 4.29 0.630 ;
        RECT 4.26 0.570 4.34 0.720 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.75 0.430 4.96 0.700 ;
        RECT 4.75 0.430 5.39 0.510 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 6.345 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 6.345 0.06 ;
    END
  END VSS

END NOR4X8

MACRO AOI21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X2 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.420 1.36 0.540 ;
        RECT 1.46 0.280 1.56 0.500 ;
        RECT 1.24 0.420 1.56 0.500 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.390 0.86 0.470 ;
        RECT 0.66 0.390 0.74 0.530 ;
        RECT 0.66 0.390 0.86 0.510 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.570 0.56 0.700 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.51 0.210 0.62 0.270 ;
        RECT 0.57 0.230 1.14 0.290 ;
        RECT 1.06 0.230 1.14 0.530 ;
        RECT 1.08 0.170 1.14 0.700 ;
        RECT 1.08 0.640 1.27 0.700 ;
        RECT 1.21 0.640 1.27 0.820 ;
    END
  END Y
END AOI21X2


MACRO NOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X2 0 0 ;
  SIZE 1.350 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.30 0.270 0.36 0.410 ;
        RECT 0.51 0.690 0.56 0.980 ;
        RECT 0.71 0.270 0.77 0.410 ;
        RECT 0.30 0.350 1.12 0.410 ;
        RECT 1.06 0.350 1.12 0.750 ;
        RECT 1.06 0.590 1.14 0.750 ;
        RECT 0.51 0.690 1.14 0.750 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.690 0.34 0.980 ;
        RECT 0.26 0.690 0.41 0.770 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.510 0.14 0.720 ;
        RECT 0.06 0.510 0.84 0.590 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.350 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.350 0.06 ;
    END
  END VSS

END NOR2X2



MACRO NOR3BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX4 0 0 ;
  SIZE 3.645 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.210 0.14 0.340 ;
        RECT 0.06 0.210 0.32 0.270 ;
        RECT 0.26 0.180 0.32 0.980 ;
        RECT 0.93 0.920 0.98 0.980 ;
        RECT 0.26 0.920 2.23 0.980 ;
        RECT 2.17 0.920 2.23 0.980 ;
        RECT 0.26 0.180 2.90 0.230 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.400 0.74 0.660 ;
        RECT 1.50 0.490 1.56 0.660 ;
        RECT 0.66 0.610 1.56 0.660 ;
        RECT 1.50 0.490 2.00 0.560 ;
        RECT 1.94 0.490 2.00 0.660 ;
        RECT 2.59 0.490 2.65 0.660 ;
        RECT 1.94 0.610 2.65 0.660 ;
        RECT 2.59 0.490 2.71 0.540 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.81 0.340 3.10 0.500 ;
        RECT 3.02 0.340 3.10 0.590 ;
        RECT 3.02 0.510 3.14 0.590 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.03 0.420 1.17 0.500 ;
        RECT 1.34 0.340 1.41 0.500 ;
        RECT 1.03 0.450 1.41 0.500 ;
        RECT 1.34 0.340 2.23 0.390 ;
        RECT 2.17 0.340 2.23 0.500 ;
        RECT 2.17 0.450 2.29 0.500 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.645 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.645 0.06 ;
    END
  END VSS

END NOR3BX4





MACRO NOR3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X4 0 0 ;
  SIZE 3.240 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.92 0.920 0.97 0.980 ;
        RECT 2.17 0.920 2.23 0.980 ;
        RECT 0.26 0.180 2.92 0.230 ;
        RECT 2.86 0.180 2.92 0.980 ;
        RECT 0.92 0.920 2.92 0.980 ;
        RECT 2.86 0.210 2.94 0.340 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.590 0.14 0.720 ;
        RECT 0.08 0.590 0.14 0.810 ;
        RECT 0.08 0.750 0.57 0.810 ;
        RECT 1.52 0.650 1.65 0.820 ;
        RECT 2.64 0.620 2.70 0.820 ;
        RECT 0.52 0.760 2.70 0.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.49 0.590 0.73 0.650 ;
        RECT 1.36 0.490 1.43 0.660 ;
        RECT 0.68 0.610 1.43 0.660 ;
        RECT 1.36 0.490 1.83 0.560 ;
        RECT 1.77 0.490 1.83 0.620 ;
        RECT 2.31 0.470 2.37 0.620 ;
        RECT 1.77 0.560 2.37 0.620 ;
        RECT 2.46 0.400 2.54 0.530 ;
        RECT 2.31 0.470 2.54 0.530 ;
        RECT 2.47 0.400 2.54 0.590 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.93 0.340 0.98 0.500 ;
        RECT 0.83 0.420 0.98 0.500 ;
        RECT 0.93 0.340 2.06 0.390 ;
        RECT 2.00 0.340 2.06 0.460 ;
        RECT 2.00 0.400 2.12 0.460 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.240 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.240 0.06 ;
    END
  END VSS

END NOR3X4

MACRO AOI31X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X4 0 0 ;
  SIZE 4.050 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.91 0.340 1.97 0.480 ;
        RECT 2.32 0.340 2.38 0.480 ;
        RECT 2.73 0.340 2.79 0.480 ;
        RECT 2.94 0.790 3.00 0.910 ;
        RECT 3.14 0.340 3.20 0.480 ;
        RECT 2.94 0.790 3.54 0.850 ;
        RECT 3.41 0.790 3.47 0.910 ;
        RECT 3.46 0.410 3.52 0.910 ;
        RECT 3.46 0.780 3.54 0.910 ;
        RECT 3.55 0.340 3.61 0.480 ;
        RECT 1.91 0.410 3.61 0.480 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.490 0.52 0.580 ;
        RECT 0.43 0.490 0.52 0.700 ;
        RECT 0.43 0.610 0.84 0.700 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.21 0.490 1.32 0.700 ;
        RECT 1.21 0.610 1.36 0.700 ;
        RECT 1.21 0.610 1.67 0.690 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.04 0.580 3.17 0.700 ;
        RECT 2.90 0.580 3.36 0.650 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.04 0.610 2.54 0.700 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.050 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.050 0.06 ;
    END
  END VSS

END AOI31X4

MACRO OAI32X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X2 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.81 0.820 0.87 0.980 ;
        RECT 1.23 0.800 1.50 0.880 ;
        RECT 0.81 0.820 1.50 0.880 ;
        RECT 1.44 0.310 1.50 0.980 ;
        RECT 1.73 0.260 1.85 0.360 ;
        RECT 1.44 0.310 2.19 0.360 ;
        RECT 2.12 0.260 2.26 0.320 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.640 0.54 0.920 ;
        RECT 0.46 0.640 0.76 0.730 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.470 1.16 0.540 ;
        RECT 0.86 0.470 0.94 0.720 ;
        RECT 0.86 0.470 1.16 0.590 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.620 1.94 0.950 ;
        RECT 1.84 0.620 2.10 0.710 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.310 0.29 0.530 ;
        RECT 0.23 0.310 1.34 0.360 ;
        RECT 1.26 0.310 1.34 0.530 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.470 1.74 0.720 ;
        RECT 1.60 0.470 2.30 0.520 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.835 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.835 0.06 ;
    END
  END VSS

END OAI32X2


MACRO NOR4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X6 0 0 ;
  SIZE 4.995 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.33 0.150 0.39 0.440 ;
        RECT 0.74 0.150 0.80 0.440 ;
        RECT 1.15 0.150 1.21 0.440 ;
        RECT 1.61 0.150 1.68 0.440 ;
        RECT 2.02 0.150 2.08 0.440 ;
        RECT 2.54 0.150 2.60 0.440 ;
        RECT 2.96 0.150 3.02 0.440 ;
        RECT 3.37 0.150 3.42 0.440 ;
        RECT 3.59 0.720 3.65 0.980 ;
        RECT 3.87 0.150 3.93 0.440 ;
        RECT 3.59 0.890 4.12 0.950 ;
        RECT 4.07 0.720 4.12 0.980 ;
        RECT 0.33 0.380 4.34 0.440 ;
        RECT 4.26 0.380 4.32 0.780 ;
        RECT 4.28 0.150 4.34 0.530 ;
        RECT 4.07 0.720 4.54 0.780 ;
        RECT 4.47 0.700 4.54 0.980 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 0.550 0.74 0.630 ;
        RECT 0.66 0.540 0.74 0.720 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.560 1.57 0.700 ;
        RECT 1.39 0.560 1.83 0.640 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.59 0.540 3.14 0.620 ;
        RECT 3.06 0.540 3.14 0.720 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.83 0.540 3.96 0.700 ;
        RECT 3.70 0.540 4.12 0.620 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.995 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.995 0.06 ;
    END
  END VSS

END NOR4X6


MACRO NAND4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X8 0 0 ;
  SIZE 6.210 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.770 0.35 0.980 ;
        RECT 0.29 0.910 0.76 0.970 ;
        RECT 0.70 0.770 0.76 0.980 ;
        RECT 1.11 0.820 1.17 0.980 ;
        RECT 1.52 0.740 1.58 0.980 ;
        RECT 1.93 0.820 1.99 0.980 ;
        RECT 0.70 0.820 2.40 0.880 ;
        RECT 2.34 0.770 2.40 0.980 ;
        RECT 2.75 0.740 2.81 0.980 ;
        RECT 2.34 0.770 3.22 0.830 ;
        RECT 3.16 0.740 3.22 0.980 ;
        RECT 3.57 0.740 3.63 0.980 ;
        RECT 3.98 0.820 4.04 0.980 ;
        RECT 4.39 0.740 4.45 0.980 ;
        RECT 4.80 0.790 4.86 0.980 ;
        RECT 3.16 0.820 5.27 0.880 ;
        RECT 5.21 0.790 5.27 0.980 ;
        RECT 5.46 0.370 5.52 0.850 ;
        RECT 5.46 0.370 5.54 0.530 ;
        RECT 5.21 0.790 5.68 0.850 ;
        RECT 5.62 0.740 5.68 0.980 ;
        RECT 4.56 0.370 5.92 0.430 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.40 0.590 1.03 0.670 ;
        RECT 0.86 0.590 0.94 0.720 ;
        RECT 0.95 0.590 1.03 0.710 ;
        RECT 0.86 0.590 1.03 0.710 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.590 1.94 0.710 ;
        RECT 1.86 0.590 2.14 0.710 ;
        RECT 2.06 0.590 2.14 0.720 ;
        RECT 1.86 0.590 2.50 0.670 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.84 0.520 3.92 0.640 ;
        RECT 3.27 0.590 3.92 0.640 ;
        RECT 3.86 0.590 3.94 0.720 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.71 0.610 5.36 0.700 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 6.210 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 6.210 0.06 ;
    END
  END VSS

END NAND4X8








MACRO NOR3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X2 0 0 ;
  SIZE 1.755 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.85 0.820 0.91 0.940 ;
        RECT 0.24 0.120 1.54 0.180 ;
        RECT 1.46 0.120 1.52 0.880 ;
        RECT 0.85 0.820 1.52 0.880 ;
        RECT 1.46 0.120 1.54 0.340 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.610 0.56 0.700 ;
        RECT 0.48 0.600 0.92 0.680 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.440 1.15 0.500 ;
        RECT 1.06 0.440 1.14 0.720 ;
        RECT 1.06 0.440 1.15 0.560 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.280 0.14 0.530 ;
        RECT 0.06 0.280 1.31 0.340 ;
        RECT 1.25 0.280 1.31 0.500 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.755 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.755 0.06 ;
    END
  END VSS

END NOR3X2





MACRO NAND4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X6 0 0 ;
  SIZE 5.130 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.720 0.49 0.980 ;
        RECT 0.84 0.700 0.90 0.980 ;
        RECT 0.43 0.890 1.31 0.950 ;
        RECT 1.25 0.700 1.31 0.980 ;
        RECT 1.80 0.820 1.86 0.980 ;
        RECT 2.29 0.700 2.34 0.980 ;
        RECT 2.69 0.720 2.75 0.980 ;
        RECT 1.25 0.820 3.23 0.880 ;
        RECT 3.17 0.750 3.23 0.980 ;
        RECT 3.17 0.750 3.63 0.810 ;
        RECT 3.58 0.700 3.63 0.980 ;
        RECT 3.83 0.320 3.88 0.440 ;
        RECT 3.58 0.890 4.12 0.950 ;
        RECT 4.07 0.720 4.12 0.980 ;
        RECT 3.83 0.380 4.32 0.440 ;
        RECT 4.26 0.320 4.32 0.880 ;
        RECT 4.26 0.590 4.34 0.720 ;
        RECT 4.07 0.820 4.54 0.880 ;
        RECT 4.47 0.700 4.54 0.980 ;
        RECT 4.68 0.150 4.74 0.460 ;
        RECT 4.26 0.400 4.74 0.460 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.540 0.74 0.620 ;
        RECT 0.66 0.540 0.74 0.760 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.540 1.74 0.720 ;
        RECT 1.66 0.570 2.06 0.650 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.73 0.540 2.92 0.620 ;
        RECT 2.86 0.570 2.94 0.720 ;
        RECT 3.02 0.530 3.10 0.650 ;
        RECT 2.83 0.570 3.10 0.650 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.73 0.610 3.96 0.700 ;
        RECT 3.86 0.540 4.16 0.620 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.130 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.130 0.06 ;
    END
  END VSS

END NAND4X6

MACRO SDFFSX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX2 0 0 ;
  SIZE 7.020 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.400 1.15 0.530 ;
        RECT 1.06 0.340 1.15 0.980 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.400 0.34 0.530 ;
        RECT 0.28 0.340 0.34 0.980 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.89 0.450 5.95 0.880 ;
        RECT 5.83 0.820 5.95 0.880 ;
        RECT 6.11 0.380 6.17 0.500 ;
        RECT 5.89 0.450 6.37 0.500 ;
        RECT 6.11 0.420 6.50 0.490 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.43 0.610 6.61 0.850 ;
        RECT 6.27 0.770 6.61 0.850 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.46 0.350 5.54 0.570 ;
        RECT 5.26 0.350 5.63 0.430 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.04 0.440 5.17 0.880 ;
        RECT 5.04 0.800 5.17 0.880 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.23 0.220 2.29 0.800 ;
        RECT 2.23 0.710 2.37 0.800 ;
        RECT 1.85 0.730 2.37 0.800 ;
        RECT 2.23 0.220 3.06 0.280 ;
        RECT 3.00 0.220 3.06 0.450 ;
        RECT 3.38 0.230 3.44 0.450 ;
        RECT 3.00 0.390 3.44 0.450 ;
        RECT 3.38 0.230 3.50 0.290 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 7.020 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 7.020 0.06 ;
    END
  END VSS

END SDFFSX2

MACRO NOR4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X4 0 0 ;
  SIZE 4.050 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.59 0.320 0.65 0.460 ;
        RECT 1.00 0.320 1.06 0.460 ;
        RECT 1.06 0.590 1.14 0.720 ;
        RECT 1.08 0.390 1.14 0.850 ;
        RECT 1.41 0.320 1.47 0.460 ;
        RECT 1.82 0.320 1.88 0.460 ;
        RECT 2.23 0.320 2.29 0.460 ;
        RECT 2.64 0.320 2.70 0.460 ;
        RECT 3.00 0.790 3.06 0.940 ;
        RECT 3.05 0.320 3.11 0.460 ;
        RECT 1.08 0.790 3.46 0.850 ;
        RECT 3.41 0.790 3.46 0.940 ;
        RECT 3.46 0.320 3.52 0.460 ;
        RECT 0.59 0.390 3.52 0.460 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.560 0.94 0.750 ;
        RECT 0.35 0.670 0.94 0.750 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.73 0.560 1.81 0.700 ;
        RECT 1.24 0.610 1.81 0.700 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.44 0.580 2.57 0.700 ;
        RECT 2.11 0.610 2.57 0.700 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.10 0.580 3.19 0.700 ;
        RECT 2.83 0.610 3.42 0.700 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.050 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.050 0.06 ;
    END
  END VSS

END NOR4X4


MACRO AOI222X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X4 0 0 ;
  SIZE 5.805 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.76 0.270 0.88 0.340 ;
        RECT 1.38 0.270 1.50 0.360 ;
        RECT 1.83 0.610 1.96 0.700 ;
        RECT 1.91 0.290 1.96 0.850 ;
        RECT 2.34 0.270 2.46 0.360 ;
        RECT 3.21 0.270 3.33 0.360 ;
        RECT 3.85 0.790 3.92 0.940 ;
        RECT 3.98 0.270 4.10 0.360 ;
        RECT 4.26 0.790 4.33 0.940 ;
        RECT 0.83 0.290 4.56 0.360 ;
        RECT 4.51 0.270 4.72 0.340 ;
        RECT 4.67 0.790 4.74 0.940 ;
        RECT 1.91 0.790 5.14 0.850 ;
        RECT 5.08 0.790 5.14 0.940 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.46 0.610 3.20 0.700 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.610 1.43 0.700 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.05 0.610 4.79 0.700 ;
    END
  END C1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.23 0.460 2.29 0.700 ;
        RECT 2.23 0.610 2.37 0.700 ;
        RECT 2.11 0.460 3.61 0.510 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.83 0.420 4.96 0.510 ;
        RECT 3.75 0.460 5.15 0.510 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.420 0.56 0.510 ;
        RECT 0.42 0.460 1.73 0.510 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.805 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.805 0.06 ;
    END
  END VSS

END AOI222X4


MACRO NOR4BBX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX2 0 0 ;
  SIZE 3.240 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.200 1.38 0.260 ;
        RECT 1.33 0.250 2.72 0.280 ;
        RECT 1.71 0.160 1.77 0.310 ;
        RECT 1.26 0.220 1.77 0.260 ;
        RECT 2.12 0.170 2.19 0.310 ;
        RECT 2.54 0.170 2.59 0.310 ;
        RECT 1.71 0.250 2.72 0.310 ;
        RECT 2.63 0.610 2.69 0.950 ;
        RECT 2.66 0.250 2.72 0.660 ;
        RECT 2.66 0.400 2.74 0.530 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.23 0.450 2.37 0.700 ;
        RECT 2.23 0.450 2.56 0.530 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.04 0.410 2.12 0.730 ;
        RECT 1.86 0.560 2.12 0.730 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.52 0.610 0.59 0.880 ;
        RECT 0.29 0.800 0.59 0.880 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.420 0.38 0.710 ;
        RECT 0.29 0.420 0.59 0.500 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.240 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.240 0.06 ;
    END
  END VSS

END NOR4BBX2




MACRO NOR4BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX2 0 0 ;
  SIZE 2.97 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.98 0.210 1.04 0.350 ;
        RECT 1.26 0.590 1.35 0.720 ;
        RECT 1.29 0.280 1.35 0.850 ;
        RECT 1.40 0.210 1.46 0.350 ;
        RECT 1.84 0.210 1.91 0.350 ;
        RECT 2.25 0.210 2.31 0.350 ;
        RECT 0.98 0.280 2.31 0.350 ;
        RECT 1.29 0.790 2.52 0.850 ;
        RECT 2.46 0.790 2.52 0.940 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.590 0.14 0.720 ;
        RECT 0.36 0.530 0.46 0.670 ;
        RECT 0.06 0.590 0.46 0.670 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.450 1.54 0.700 ;
        RECT 1.64 0.600 1.77 0.700 ;
        RECT 1.46 0.610 1.77 0.700 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.87 0.450 2.04 0.700 ;
        RECT 1.87 0.610 2.20 0.700 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.30 0.450 2.47 0.700 ;
        RECT 2.30 0.610 2.56 0.700 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.97 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.97 0.06 ;
    END
  END VSS

END NOR4BX2


MACRO NAND4BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX2 0 0 ;
  SIZE 2.97 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.89 0.910 0.94 0.980 ;
        RECT 1.18 0.460 1.24 0.980 ;
        RECT 1.26 0.910 1.35 0.980 ;
        RECT 1.29 0.910 1.35 0.980 ;
        RECT 1.71 0.910 1.77 0.980 ;
        RECT 0.89 0.910 2.21 0.980 ;
        RECT 2.12 0.910 2.21 0.980 ;
        RECT 2.22 0.260 2.28 0.510 ;
        RECT 1.18 0.460 2.28 0.510 ;
        RECT 2.22 0.260 2.35 0.320 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.04 0.500 0.26 0.590 ;
        RECT 0.18 0.500 0.26 0.700 ;
        RECT 0.18 0.610 0.42 0.700 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.34 0.610 1.56 0.810 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.67 0.610 1.96 0.810 ;
        RECT 1.67 0.650 2.04 0.810 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.16 0.610 2.57 0.770 ;
        RECT 2.15 0.690 2.57 0.770 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.97 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.97 0.06 ;
    END
  END VSS

END NAND4BX2

MACRO NAND4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X4 0 0 ;
  SIZE 4.185 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.770 0.34 0.980 ;
        RECT 0.69 0.770 0.76 0.980 ;
        RECT 1.08 0.460 1.14 0.910 ;
        RECT 1.06 0.790 1.19 0.910 ;
        RECT 0.28 0.770 1.14 0.830 ;
        RECT 1.13 0.790 1.19 0.980 ;
        RECT 1.54 0.790 1.60 0.980 ;
        RECT 1.98 0.790 2.04 0.980 ;
        RECT 2.40 0.790 2.46 0.980 ;
        RECT 2.75 0.330 2.81 0.510 ;
        RECT 1.08 0.460 2.81 0.510 ;
        RECT 2.97 0.790 3.03 0.980 ;
        RECT 3.21 0.250 3.27 0.380 ;
        RECT 1.06 0.790 3.44 0.850 ;
        RECT 3.38 0.790 3.44 0.980 ;
        RECT 3.63 0.250 3.69 0.380 ;
        RECT 2.75 0.330 3.69 0.380 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.420 0.73 0.500 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.610 1.74 0.700 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.83 0.610 2.96 0.700 ;
        RECT 2.91 0.490 2.96 0.700 ;
        RECT 2.10 0.630 2.96 0.700 ;
        RECT 2.91 0.490 3.02 0.540 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 0.490 3.54 0.700 ;
        RECT 3.10 0.610 3.54 0.700 ;
        RECT 3.46 0.490 3.58 0.570 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.185 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.185 0.06 ;
    END
  END VSS

END NAND4X4





MACRO TLATNTSCAX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX3 0 0 ;
  SIZE 4.185 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.42 0.700 3.48 0.980 ;
        RECT 3.46 0.320 3.52 0.760 ;
        RECT 3.46 0.400 3.54 0.530 ;
        RECT 3.42 0.700 3.88 0.760 ;
        RECT 3.83 0.700 3.88 0.980 ;
        RECT 3.87 0.320 3.93 0.460 ;
        RECT 3.46 0.400 3.93 0.460 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.250 0.77 0.730 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.400 0.52 0.730 ;
        RECT 0.46 0.250 0.54 0.530 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.330 0.17 0.700 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.185 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.185 0.06 ;
    END
  END VSS

END TLATNTSCAX3






















MACRO OAI33X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X2 0 0 ;
  SIZE 4.590 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.03 0.800 3.17 0.880 ;
        RECT 3.97 0.740 4.03 0.860 ;
        RECT 2.84 0.800 4.03 0.860 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 0.790 2.23 0.850 ;
        RECT 2.04 0.790 2.23 0.880 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 0.640 2.74 0.910 ;
        RECT 2.66 0.780 2.74 0.910 ;
        RECT 2.68 0.640 3.87 0.710 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.610 1.94 0.680 ;
        RECT 1.64 0.610 1.94 0.700 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.46 0.490 2.54 0.720 ;
        RECT 2.46 0.490 3.71 0.540 ;
    END
  END B2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.420 0.56 0.500 ;
        RECT 0.33 0.450 1.50 0.500 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.48 0.210 2.59 0.320 ;
        RECT 0.64 0.230 2.59 0.320 ;
        RECT 2.54 0.210 2.59 0.380 ;
        RECT 2.92 0.210 3.04 0.380 ;
        RECT 3.35 0.210 3.48 0.380 ;
        RECT 3.79 0.210 3.87 0.380 ;
        RECT 2.54 0.330 3.87 0.380 ;
        RECT 3.79 0.210 3.92 0.270 ;
        RECT 4.13 0.370 4.19 0.980 ;
        RECT 4.19 0.250 4.25 0.440 ;
        RECT 3.81 0.370 4.25 0.440 ;
        RECT 4.24 0.190 4.29 0.310 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.590 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.590 0.06 ;
    END
  END VSS

END OAI33X2






















MACRO SEDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX4 0 0 ;
  SIZE 8.370 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.07 0.450 7.13 0.690 ;
        RECT 7.01 0.630 7.13 0.690 ;
        RECT 7.63 0.420 7.97 0.500 ;
        RECT 7.07 0.450 7.97 0.500 ;
        RECT 7.91 0.420 7.97 0.540 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.39 0.610 7.56 0.760 ;
        RECT 7.39 0.610 7.81 0.690 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.42 0.490 6.50 0.740 ;
        RECT 6.42 0.610 6.75 0.740 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.510 5.34 0.980 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.83 0.580 5.16 0.700 ;
        RECT 5.08 0.510 5.16 0.760 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.340 0.34 0.980 ;
        RECT 0.26 0.400 0.34 0.530 ;
        RECT 0.26 0.470 0.74 0.530 ;
        RECT 0.69 0.340 0.74 0.980 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 8.370 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 8.370 0.06 ;
    END
  END VSS

END SEDFFHQX4
















MACRO AOI32X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X2 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.50 0.230 1.56 0.880 ;
        RECT 1.44 0.800 1.56 0.880 ;
        RECT 1.44 0.800 1.79 0.860 ;
        RECT 1.73 0.800 1.79 0.980 ;
        RECT 0.81 0.230 2.02 0.290 ;
        RECT 1.73 0.900 2.20 0.970 ;
        RECT 2.14 0.900 2.20 0.980 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.52 0.720 0.60 0.880 ;
        RECT 0.43 0.800 0.60 0.880 ;
        RECT 0.52 0.720 0.85 0.790 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.52 0.560 1.14 0.610 ;
        RECT 1.06 0.560 1.14 0.720 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.89 0.680 2.34 0.800 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.390 0.42 0.620 ;
        RECT 0.36 0.390 1.34 0.460 ;
        RECT 1.26 0.390 1.34 0.620 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.67 0.420 1.79 0.600 ;
        RECT 1.67 0.420 2.54 0.500 ;
        RECT 2.42 0.420 2.54 0.600 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.835 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.835 0.06 ;
    END
  END VSS

END AOI32X2


MACRO OR3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X4 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.91 0.710 0.96 0.980 ;
        RECT 0.92 0.200 1.03 0.260 ;
        RECT 0.98 0.220 1.49 0.280 ;
        RECT 1.31 0.870 1.38 0.980 ;
        RECT 0.91 0.710 1.49 0.770 ;
        RECT 1.37 0.160 1.43 0.280 ;
        RECT 1.43 0.220 1.49 0.930 ;
        RECT 1.31 0.870 1.49 0.930 ;
        RECT 1.43 0.400 1.74 0.460 ;
        RECT 1.66 0.400 1.74 0.530 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.540 0.74 0.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.780 0.34 0.910 ;
        RECT 0.32 0.470 0.40 0.860 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.410 0.14 0.910 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS

END OR3X4

























MACRO TLATNTSCAX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX8 0 0 ;
  SIZE 5.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.760 3.74 0.910 ;
        RECT 3.68 0.320 3.74 0.980 ;
        RECT 4.09 0.760 4.15 0.980 ;
        RECT 4.06 0.350 4.18 0.400 ;
        RECT 4.50 0.760 4.56 0.980 ;
        RECT 4.47 0.350 4.59 0.420 ;
        RECT 4.13 0.360 4.97 0.420 ;
        RECT 3.66 0.760 4.97 0.820 ;
        RECT 4.91 0.300 4.97 0.980 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.250 0.74 0.530 ;
        RECT 0.68 0.400 0.76 0.740 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 0.250 0.53 0.740 ;
        RECT 0.45 0.250 0.54 0.530 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.270 0.18 0.700 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.400 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.400 0.06 ;
    END
  END VSS

END TLATNTSCAX8






















MACRO AOI222X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X2 0 0 ;
  SIZE 3.375 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.590 1.34 0.720 ;
        RECT 1.28 0.250 1.34 0.860 ;
        RECT 1.28 0.800 2.50 0.860 ;
        RECT 2.44 0.800 2.50 0.960 ;
        RECT 0.70 0.250 2.67 0.310 ;
        RECT 2.44 0.820 2.91 0.880 ;
        RECT 2.85 0.810 2.91 0.940 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 0.610 2.13 0.700 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.620 0.83 0.750 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.56 0.590 2.73 0.720 ;
        RECT 2.56 0.610 2.74 0.700 ;
    END
  END C1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.420 0.56 0.540 ;
        RECT 0.51 0.410 0.95 0.490 ;
        RECT 0.86 0.440 1.06 0.510 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.83 0.420 1.96 0.510 ;
        RECT 1.50 0.440 2.13 0.510 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.23 0.420 2.40 0.510 ;
        RECT 2.23 0.420 2.90 0.490 ;
        RECT 2.84 0.480 3.02 0.540 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.375 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.375 0.06 ;
    END
  END VSS

END AOI222X2







MACRO NAND2BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX4 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.250 0.14 0.980 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.420 0.47 0.800 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.85 0.380 1.94 0.730 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS

END NAND2BX4


MACRO AOI33X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X2 0 0 ;
  SIZE 3.240 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.50 0.140 1.56 0.880 ;
        RECT 1.44 0.800 1.56 0.880 ;
        RECT 1.44 0.820 1.79 0.880 ;
        RECT 1.73 0.820 1.79 0.970 ;
        RECT 0.76 0.140 2.19 0.200 ;
        RECT 2.16 0.840 2.22 0.970 ;
        RECT 1.73 0.840 2.65 0.900 ;
        RECT 2.59 0.840 2.65 0.970 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.69 0.610 0.96 0.720 ;
        RECT 0.69 0.610 1.16 0.700 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.90 0.610 2.14 0.730 ;
        RECT 1.90 0.610 2.36 0.700 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 0.460 2.54 0.510 ;
        RECT 2.46 0.460 2.54 0.720 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.460 0.54 0.720 ;
        RECT 0.42 0.460 1.11 0.510 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.290 0.32 0.520 ;
        RECT 0.26 0.290 1.32 0.360 ;
        RECT 1.26 0.290 1.32 0.530 ;
        RECT 1.26 0.400 1.34 0.530 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.68 0.290 1.74 0.530 ;
        RECT 1.66 0.400 1.74 0.530 ;
        RECT 1.68 0.290 2.70 0.360 ;
        RECT 2.64 0.290 2.70 0.530 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.240 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.240 0.06 ;
    END
  END VSS

END AOI33X2















MACRO TLATNTSCAX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX6 0 0 ;
  SIZE 5.130 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.150 3.92 0.980 ;
        RECT 3.86 0.560 3.94 0.720 ;
        RECT 4.27 0.150 4.33 0.980 ;
        RECT 3.86 0.560 4.74 0.620 ;
        RECT 4.63 0.400 4.70 0.620 ;
        RECT 4.68 0.150 4.74 0.460 ;
        RECT 4.68 0.560 4.74 0.980 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.250 0.74 0.750 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.250 0.54 0.750 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.280 0.20 0.700 ;
#        RECT 0.035 0.815 0.2 0.895 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.130 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.130 0.06 ;
    END
  END VSS

END TLATNTSCAX6















MACRO OAI211X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X2 0 0 ;
  SIZE 2.565 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.860 0.70 0.980 ;
        RECT 1.28 0.440 1.34 0.920 ;
        RECT 1.26 0.780 1.34 0.920 ;
        RECT 1.34 0.860 1.40 0.980 ;
        RECT 0.64 0.860 1.81 0.920 ;
        RECT 1.75 0.860 1.81 0.980 ;
        RECT 1.96 0.260 2.02 0.490 ;
        RECT 1.28 0.440 2.02 0.490 ;
        RECT 1.96 0.260 2.13 0.320 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.610 0.54 0.910 ;
        RECT 0.46 0.610 0.74 0.700 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.590 0.34 0.720 ;
        RECT 0.28 0.440 0.36 0.680 ;
        RECT 0.28 0.440 0.97 0.510 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.600 1.85 0.760 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.12 0.410 2.19 0.700 ;
        RECT 2.12 0.590 2.34 0.700 ;
        RECT 2.26 0.590 2.34 0.770 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.565 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.565 0.06 ;
    END
  END VSS

END OAI211X2































MACRO SEDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX8 0 0 ;
  SIZE 8.910 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.76 0.440 7.82 0.810 ;
        RECT 8.04 0.420 8.16 0.500 ;
        RECT 7.76 0.440 8.16 0.490 ;
        RECT 8.04 0.450 8.61 0.500 ;
        RECT 8.55 0.450 8.61 0.570 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.14 0.610 8.45 0.700 ;
        RECT 8.37 0.610 8.45 0.870 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.420 7.34 0.920 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.08 0.440 6.17 0.750 ;
        RECT 6.04 0.610 6.17 0.750 ;
        RECT 6.08 0.440 6.30 0.520 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.58 0.500 2.74 0.720 ;
        RECT 2.66 0.500 2.74 0.920 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.400 0.14 0.530 ;
        RECT 0.08 0.340 0.14 0.980 ;
        RECT 0.06 0.450 0.55 0.500 ;
        RECT 0.49 0.340 0.55 0.980 ;
        RECT 0.90 0.340 0.96 0.980 ;
        RECT 0.49 0.540 1.32 0.600 ;
        RECT 1.27 0.380 1.32 0.760 ;
        RECT 1.31 0.330 1.37 0.450 ;
        RECT 1.31 0.700 1.37 0.980 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 8.910 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 8.910 0.06 ;
    END
  END VSS

END SEDFFHQX8


MACRO TLATNTSCAX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX4 0 0 ;
  SIZE 4.320 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 0.800 0.81 0.980 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.610 0.93 0.710 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.780 0.14 0.950 ;
        RECT 0.10 0.490 0.17 0.860 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.44 0.270 3.52 0.380 ;
        RECT 3.44 0.770 3.50 0.980 ;
        RECT 3.46 0.270 3.52 0.530 ;
        RECT 3.46 0.400 3.54 0.530 ;
        RECT 3.49 0.470 3.55 0.830 ;
        RECT 3.46 0.470 3.92 0.530 ;
        RECT 3.85 0.270 3.92 0.980 ;
    END
  END ECK
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.320 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.320 0.06 ;
    END
  END VSS

END TLATNTSCAX4








MACRO OR4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X2 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.200 1.74 0.980 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.400 0.74 0.530 ;
        RECT 0.66 0.400 0.92 0.480 ;
        RECT 0.84 0.280 0.92 0.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.280 0.56 0.760 ;
        RECT 0.46 0.590 0.56 0.760 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.280 0.36 0.760 ;
        RECT 0.26 0.590 0.36 0.760 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.20 0.150 1.27 0.560 ;
        RECT 1.20 0.420 1.36 0.500 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS

END OR4X2














MACRO AOI221X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X4 0 0 ;
  SIZE 4.725 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.76 0.250 0.88 0.310 ;
        RECT 1.38 0.250 1.50 0.330 ;
        RECT 1.83 0.420 1.96 0.500 ;
        RECT 1.91 0.270 1.96 0.850 ;
        RECT 2.37 0.250 2.49 0.330 ;
        RECT 3.13 0.250 3.25 0.330 ;
        RECT 3.67 0.250 3.79 0.330 ;
        RECT 3.83 0.790 3.90 0.940 ;
        RECT 0.83 0.270 4.17 0.330 ;
        RECT 4.12 0.250 4.24 0.310 ;
        RECT 1.91 0.790 4.30 0.850 ;
        RECT 4.25 0.790 4.30 0.940 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.69 0.610 1.43 0.700 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.50 0.610 3.18 0.700 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.420 0.36 0.500 ;
        RECT 0.23 0.450 1.73 0.500 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.42 0.460 3.48 0.700 ;
        RECT 2.09 0.460 3.54 0.510 ;
        RECT 3.42 0.610 3.56 0.700 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.83 0.420 3.96 0.700 ;
        RECT 3.83 0.430 4.20 0.510 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.725 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.725 0.06 ;
    END
  END VSS

END AOI221X4












MACRO NAND3BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX4 0 0 ;
  SIZE 3.240 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.210 0.14 0.340 ;
        RECT 0.08 0.210 0.14 0.890 ;
        RECT 0.08 0.830 0.36 0.890 ;
        RECT 0.30 0.830 0.36 0.980 ;
        RECT 0.71 0.920 0.77 0.980 ;
        RECT 1.12 0.920 1.18 0.980 ;
        RECT 1.53 0.920 1.59 0.980 ;
        RECT 0.06 0.210 1.95 0.270 ;
        RECT 1.94 0.920 2.00 0.980 ;
        RECT 0.30 0.920 2.41 0.980 ;
        RECT 2.35 0.920 2.41 0.980 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.420 0.56 0.510 ;
        RECT 0.40 0.460 0.72 0.510 ;
        RECT 0.66 0.460 0.72 0.660 ;
        RECT 0.66 0.610 1.28 0.660 ;
        RECT 1.23 0.540 1.67 0.610 ;
        RECT 1.60 0.610 2.27 0.660 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.37 0.420 2.56 0.500 ;
        RECT 2.48 0.420 2.56 0.600 ;
        RECT 2.48 0.510 2.77 0.600 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.83 0.420 0.96 0.500 ;
        RECT 0.82 0.450 1.12 0.500 ;
        RECT 1.06 0.380 1.82 0.450 ;
        RECT 1.77 0.450 1.89 0.500 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.240 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.240 0.06 ;
    END
  END VSS

END NAND3BX4

















MACRO TLATNTSCAX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX2 0 0 ;
  SIZE 4.050 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.210 3.34 0.980 ;
        RECT 3.26 0.210 3.36 0.330 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.250 0.74 0.750 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.250 0.54 0.750 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.10 0.310 0.20 0.750 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.050 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.050 0.06 ;
    END
  END VSS

END TLATNTSCAX2





MACRO SEDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX2 0 0 ;
  SIZE 7.155 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.290 3.14 0.820 ;
        RECT 3.06 0.290 3.19 0.370 ;
        RECT 3.06 0.740 3.27 0.820 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.48 0.470 6.56 0.760 ;
        RECT 6.48 0.590 6.77 0.760 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.500 2.96 0.720 ;
        RECT 2.88 0.500 2.96 0.980 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.62 0.420 1.77 0.700 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.380 0.74 0.880 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.420 0.36 0.500 ;
        RECT 0.50 0.220 0.56 0.490 ;
        RECT 0.23 0.420 0.56 0.490 ;
        RECT 0.50 0.220 0.96 0.280 ;
        RECT 0.90 0.220 0.96 0.460 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 7.155 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 7.155 0.06 ;
    END
  END VSS

END SEDFFHQX2


















MACRO TLATNTSCAX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX20 0 0 ;
  SIZE 8.910 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.150 5.32 0.980 ;
        RECT 5.26 0.560 5.34 0.980 ;
        RECT 5.67 0.150 5.73 0.980 ;
        RECT 6.04 0.400 6.09 0.620 ;
        RECT 6.08 0.150 6.14 0.460 ;
        RECT 6.08 0.560 6.14 0.980 ;
        RECT 6.49 0.150 6.55 0.980 ;
        RECT 6.90 0.150 6.96 0.980 ;
        RECT 7.31 0.150 7.37 0.980 ;
        RECT 7.72 0.150 7.78 0.980 ;
        RECT 8.13 0.150 8.19 0.980 ;
        RECT 5.26 0.560 8.60 0.620 ;
        RECT 8.49 0.400 8.55 0.620 ;
        RECT 8.54 0.150 8.60 0.460 ;
        RECT 8.54 0.560 8.60 0.980 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.74 0.470 0.96 0.700 ;
        RECT 0.69 0.610 1.05 0.700 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.590 0.54 0.750 ;
        RECT 0.52 0.310 0.59 0.670 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.780 0.14 0.940 ;
        RECT 0.12 0.500 0.20 0.860 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 8.910 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 8.910 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal2 ;
        RECT 2.51 0.225 2.61 0.975 ;
        RECT 3.20 0.225 3.32 0.775 ;
        RECT 4.71 0.225 4.81 0.975 ;
        RECT 5.71 0.325 5.81 0.875 ;
        RECT 1.42 0.325 1.52 0.875 ;
  END
END TLATNTSCAX20


MACRO AOI211X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X2 0 0 ;
  SIZE 2.160 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 0.250 0.67 0.310 ;
        RECT 1.06 0.270 1.14 0.530 ;
        RECT 1.08 0.270 1.14 0.800 ;
        RECT 1.20 0.250 1.31 0.330 ;
        RECT 1.08 0.740 1.73 0.800 ;
        RECT 0.62 0.270 1.69 0.330 ;
        RECT 1.67 0.740 1.73 0.980 ;
        RECT 1.64 0.250 1.75 0.310 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.53 0.610 0.90 0.720 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.420 0.91 0.500 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.420 1.60 0.500 ;
        RECT 1.44 0.420 1.60 0.640 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.70 0.420 1.94 0.600 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.160 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.160 0.06 ;
    END
  END VSS

END AOI211X2



MACRO NAND2BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX2 0 0 ;
  SIZE 1.350 BY 1.2 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.350 0.15 0.980 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.03 0.480 1.11 0.980 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.460 0.56 0.980 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 1.350 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 1.350 0.06 ;
    END
  END VSS

END NAND2BX2










MACRO OAI21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X4 0 0 ;
  SIZE 2.97 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.63 0.820 0.69 0.980 ;
        RECT 1.25 0.820 1.31 0.980 ;
        RECT 1.86 0.820 1.92 0.980 ;
        RECT 1.88 0.270 1.94 0.980 ;
        RECT 0.63 0.820 1.94 0.880 ;
        RECT 1.86 0.830 1.94 0.980 ;
        RECT 1.88 0.270 2.05 0.380 ;
        RECT 1.86 0.830 2.33 0.890 ;
        RECT 2.27 0.830 2.33 0.980 ;
        RECT 1.88 0.330 2.38 0.380 ;
        RECT 2.33 0.270 2.46 0.340 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.610 0.68 0.710 ;
        RECT 0.43 0.630 1.27 0.710 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.21 0.460 0.34 0.520 ;
        RECT 0.83 0.460 0.95 0.530 ;
        RECT 0.30 0.460 1.64 0.510 ;
        RECT 1.57 0.460 1.64 0.650 ;
        RECT 1.57 0.590 1.74 0.650 ;
        RECT 1.66 0.590 1.74 0.720 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.04 0.490 2.12 0.740 ;
        RECT 2.04 0.610 2.37 0.700 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.97 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.97 0.06 ;
    END
  END VSS

END OAI21X4


MACRO NAND4BBX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX2 0 0 ;
  SIZE 3.375 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 0.800 1.61 0.980 ;
        RECT 1.55 0.800 1.77 0.960 ;
        RECT 1.96 0.890 2.02 0.980 ;
        RECT 2.37 0.890 2.43 0.980 ;
        RECT 2.82 0.890 2.88 0.980 ;
        RECT 2.87 0.240 2.92 0.960 ;
        RECT 1.55 0.890 2.92 0.960 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.320 2.74 0.530 ;
        RECT 2.69 0.450 2.77 0.790 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 0.500 2.33 0.790 ;
        RECT 2.25 0.590 2.54 0.790 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.56 0.610 0.65 0.970 ;
        RECT 0.56 0.800 0.80 0.970 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.610 0.47 0.700 ;
        RECT 0.39 0.610 0.47 0.970 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 3.375 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 3.375 0.06 ;
    END
  END VSS

END NAND4BBX2





MACRO OAI21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X2 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.940 0.70 0.980 ;
        RECT 1.06 0.590 1.14 0.720 ;
        RECT 1.06 0.660 1.30 0.720 ;
        RECT 1.20 0.940 1.25 0.980 ;
        RECT 1.24 0.400 1.30 0.980 ;
        RECT 0.65 0.940 1.30 0.980 ;
        RECT 1.32 0.340 1.39 0.460 ;
        RECT 1.24 0.400 1.39 0.460 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.760 0.54 0.980 ;
        RECT 0.46 0.760 0.70 0.840 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 0.580 0.94 0.660 ;
        RECT 0.86 0.580 0.94 0.720 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.40 0.560 1.48 0.980 ;
        RECT 1.40 0.590 1.54 0.720 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.025 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.025 0.06 ;
    END
  END VSS

END OAI21X2

MACRO NAND4BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX4 0 0 ;
  SIZE 4.590 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.69 0.760 0.74 0.980 ;
        RECT 1.09 0.760 1.16 0.980 ;
        RECT 1.48 0.460 1.54 0.910 ;
        RECT 1.46 0.790 1.58 0.910 ;
        RECT 0.69 0.760 1.54 0.820 ;
        RECT 1.52 0.790 1.58 0.980 ;
        RECT 1.93 0.790 1.99 0.980 ;
        RECT 2.34 0.790 2.40 0.980 ;
        RECT 2.75 0.790 2.81 0.980 ;
        RECT 3.10 0.310 3.16 0.510 ;
        RECT 1.48 0.460 3.16 0.510 ;
        RECT 3.31 0.790 3.37 0.980 ;
        RECT 3.54 0.220 3.59 0.360 ;
        RECT 1.46 0.790 3.77 0.850 ;
        RECT 3.71 0.790 3.77 0.980 ;
        RECT 3.97 0.220 4.03 0.360 ;
        RECT 3.10 0.310 4.03 0.360 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.400 0.14 0.530 ;
        RECT 0.10 0.450 0.18 0.860 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 0.610 2.14 0.700 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.04 0.610 3.32 0.700 ;
        RECT 3.26 0.470 3.32 0.700 ;
        RECT 2.45 0.630 3.32 0.700 ;
        RECT 3.26 0.470 3.38 0.520 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.62 0.470 3.77 0.700 ;
        RECT 3.44 0.610 3.77 0.700 ;
        RECT 3.62 0.470 3.92 0.540 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 4.590 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 4.590 0.06 ;
    END
  END VSS

END NAND4BX4



MACRO OA21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X4 0 0 ;
  SIZE 2.430 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.20 0.740 1.26 0.980 ;
        RECT 1.30 0.340 1.36 0.480 ;
        RECT 1.61 0.740 1.67 0.980 ;
        RECT 1.30 0.420 1.81 0.480 ;
        RECT 1.71 0.340 1.77 0.480 ;
        RECT 1.75 0.420 1.81 0.800 ;
        RECT 1.75 0.590 1.94 0.800 ;
        RECT 1.20 0.740 1.94 0.800 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.430 0.14 0.930 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.430 0.60 0.510 ;
        RECT 0.43 0.430 0.60 0.700 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.72 0.410 0.80 0.670 ;
        RECT 0.72 0.590 0.94 0.670 ;
        RECT 0.86 0.590 0.94 0.770 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 2.430 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 2.430 0.06 ;
    END
  END VSS

END OA21X4




MACRO TLATNTSCAX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX12 0 0 ;
  SIZE 6.615 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.24 0.150 4.29 0.460 ;
        RECT 4.24 0.670 4.29 0.980 ;
        RECT 4.24 0.670 4.30 0.730 ;
        RECT 4.26 0.400 4.32 0.720 ;
        RECT 4.26 0.590 4.34 0.720 ;
        RECT 4.64 0.150 4.71 0.980 ;
        RECT 5.05 0.150 5.12 0.980 ;
        RECT 5.46 0.150 5.53 0.980 ;
        RECT 5.83 0.590 5.89 0.810 ;
        RECT 5.88 0.150 5.94 0.650 ;
        RECT 4.26 0.590 5.94 0.650 ;
        RECT 5.88 0.750 5.94 0.980 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.250 0.74 0.530 ;
        RECT 0.67 0.250 0.74 0.740 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.250 0.54 0.740 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.280 0.14 0.700 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 6.615 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 6.615 0.06 ;
    END
  END VSS
  OBS
      LAYER Metal2 ;
        RECT 2.51 0.225 2.61 0.975 ;
        RECT 3.20 0.225 3.32 0.775 ;
        RECT 4.71 0.225 4.81 0.975 ;
        RECT 5.71 0.325 5.81 0.875 ;
        RECT 1.42 0.325 1.52 0.875 ;
  END
END TLATNTSCAX12




MACRO SDFFRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX2 0 0 ;
  SIZE 5.94 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.220 0.34 0.800 ;
        RECT 0.26 0.730 0.34 0.980 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.78 0.450 4.84 0.720 ;
        RECT 5.04 0.420 5.17 0.500 ;
        RECT 4.78 0.450 5.20 0.500 ;
        RECT 5.14 0.460 5.47 0.510 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.20 0.610 5.61 0.730 ;
        RECT 5.14 0.640 5.61 0.730 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.400 4.34 0.530 ;
        RECT 4.26 0.400 4.52 0.480 ;
        RECT 4.44 0.400 4.52 0.670 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.48 0.590 1.67 0.790 ;
        RECT 1.48 0.610 1.85 0.790 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.59 0.460 0.74 0.720 ;
        RECT 0.66 0.460 0.74 0.890 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 1.14 5.94 1.2 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
	RECT 0.00 0.00 5.94 0.06 ;
    END
  END VSS

END SDFFRHQX2



MACRO MEM1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM1 0 0 ;
  SIZE 426.965 BY 114.215 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 77.64 12.66 78.30 ;
      LAYER Metal6 ;
        RECT 12.00 77.64 12.66 78.30 ;
      LAYER Metal3 ;
        RECT 12.00 77.64 12.66 78.30 ;
      LAYER Metal4 ;
        RECT 12.00 77.64 12.66 78.30 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 71.52 12.66 72.18 ;
      LAYER Metal6 ;
        RECT 12.00 71.52 12.66 72.18 ;
      LAYER Metal3 ;
        RECT 12.00 71.52 12.66 72.18 ;
      LAYER Metal4 ;
        RECT 12.00 71.52 12.66 72.18 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 68.42 12.66 69.08 ;
      LAYER Metal6 ;
        RECT 12.00 68.42 12.66 69.08 ;
      LAYER Metal3 ;
        RECT 12.00 68.42 12.66 69.08 ;
      LAYER Metal4 ;
        RECT 12.00 68.42 12.66 69.08 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 62.30 12.66 62.96 ;
      LAYER Metal6 ;
        RECT 12.00 62.30 12.66 62.96 ;
      LAYER Metal3 ;
        RECT 12.00 62.30 12.66 62.96 ;
      LAYER Metal4 ;
        RECT 12.00 62.30 12.66 62.96 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 59.28 12.66 59.94 ;
      LAYER Metal6 ;
        RECT 12.00 59.28 12.66 59.94 ;
      LAYER Metal3 ;
        RECT 12.00 59.28 12.66 59.94 ;
      LAYER Metal4 ;
        RECT 12.00 59.28 12.66 59.94 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 56.18 12.66 56.84 ;
      LAYER Metal6 ;
        RECT 12.00 56.18 12.66 56.84 ;
      LAYER Metal3 ;
        RECT 12.00 56.18 12.66 56.84 ;
      LAYER Metal4 ;
        RECT 12.00 56.18 12.66 56.84 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 50.06 12.66 50.72 ;
      LAYER Metal6 ;
        RECT 12.00 50.06 12.66 50.72 ;
      LAYER Metal3 ;
        RECT 12.00 50.06 12.66 50.72 ;
      LAYER Metal4 ;
        RECT 12.00 50.06 12.66 50.72 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 47.04 12.66 47.70 ;
      LAYER Metal6 ;
        RECT 12.00 47.04 12.66 47.70 ;
      LAYER Metal3 ;
        RECT 12.00 47.04 12.66 47.70 ;
      LAYER Metal4 ;
        RECT 12.00 47.04 12.66 47.70 ;
    END
  END A[7]
  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 228.44 12.00 229.09 12.66 ;
      LAYER Metal6 ;
        RECT 228.44 12.00 229.09 12.66 ;
      LAYER Metal3 ;
        RECT 228.44 12.00 229.09 12.66 ;
      LAYER Metal4 ;
        RECT 228.44 12.00 229.09 12.66 ;
    END
  END CE
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal5 ;
        RECT 238.18 12.00 238.84 12.66 ;
      LAYER Metal6 ;
        RECT 238.18 12.00 238.84 12.66 ;
      LAYER Metal3 ;
        RECT 238.18 12.00 238.84 12.66 ;
      LAYER Metal4 ;
        RECT 238.18 12.00 238.84 12.66 ;
    END
  END CK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 20.48 12.00 21.14 12.66 ;
      LAYER Metal6 ;
        RECT 20.48 12.00 21.14 12.66 ;
      LAYER Metal3 ;
        RECT 20.48 12.00 21.14 12.66 ;
      LAYER Metal4 ;
        RECT 20.48 12.00 21.14 12.66 ;
    END
  END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 129.00 12.00 129.66 12.66 ;
      LAYER Metal6 ;
        RECT 129.00 12.00 129.66 12.66 ;
      LAYER Metal3 ;
        RECT 129.00 12.00 129.66 12.66 ;
      LAYER Metal4 ;
        RECT 129.00 12.00 129.66 12.66 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 137.04 12.00 137.70 12.66 ;
      LAYER Metal6 ;
        RECT 137.04 12.00 137.70 12.66 ;
      LAYER Metal3 ;
        RECT 137.04 12.00 137.70 12.66 ;
      LAYER Metal4 ;
        RECT 137.04 12.00 137.70 12.66 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 151.34 12.00 152.00 12.66 ;
      LAYER Metal6 ;
        RECT 151.34 12.00 152.00 12.66 ;
      LAYER Metal3 ;
        RECT 151.34 12.00 152.00 12.66 ;
      LAYER Metal4 ;
        RECT 151.34 12.00 152.00 12.66 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 159.38 12.00 160.04 12.66 ;
      LAYER Metal6 ;
        RECT 159.38 12.00 160.04 12.66 ;
      LAYER Metal3 ;
        RECT 159.38 12.00 160.04 12.66 ;
      LAYER Metal4 ;
        RECT 159.38 12.00 160.04 12.66 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 172.62 12.00 173.28 12.66 ;
      LAYER Metal6 ;
        RECT 172.62 12.00 173.28 12.66 ;
      LAYER Metal3 ;
        RECT 172.62 12.00 173.28 12.66 ;
      LAYER Metal4 ;
        RECT 172.62 12.00 173.28 12.66 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 180.66 12.00 181.32 12.66 ;
      LAYER Metal6 ;
        RECT 180.66 12.00 181.32 12.66 ;
      LAYER Metal3 ;
        RECT 180.66 12.00 181.32 12.66 ;
      LAYER Metal4 ;
        RECT 180.66 12.00 181.32 12.66 ;
    END
  END D[15]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 245.65 12.00 246.31 12.66 ;
      LAYER Metal6 ;
        RECT 245.65 12.00 246.31 12.66 ;
      LAYER Metal3 ;
        RECT 245.65 12.00 246.31 12.66 ;
      LAYER Metal4 ;
        RECT 245.65 12.00 246.31 12.66 ;
    END
  END D[16]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 253.69 12.00 254.34 12.66 ;
      LAYER Metal6 ;
        RECT 253.69 12.00 254.34 12.66 ;
      LAYER Metal3 ;
        RECT 253.69 12.00 254.34 12.66 ;
      LAYER Metal4 ;
        RECT 253.69 12.00 254.34 12.66 ;
    END
  END D[17]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 266.93 12.00 267.58 12.66 ;
      LAYER Metal6 ;
        RECT 266.93 12.00 267.58 12.66 ;
      LAYER Metal3 ;
        RECT 266.93 12.00 267.58 12.66 ;
      LAYER Metal4 ;
        RECT 266.93 12.00 267.58 12.66 ;
    END
  END D[18]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 274.96 12.00 275.62 12.66 ;
      LAYER Metal6 ;
        RECT 274.96 12.00 275.62 12.66 ;
      LAYER Metal3 ;
        RECT 274.96 12.00 275.62 12.66 ;
      LAYER Metal4 ;
        RECT 274.96 12.00 275.62 12.66 ;
    END
  END D[19]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 28.52 12.00 29.18 12.66 ;
      LAYER Metal6 ;
        RECT 28.52 12.00 29.18 12.66 ;
      LAYER Metal3 ;
        RECT 28.52 12.00 29.18 12.66 ;
      LAYER Metal4 ;
        RECT 28.52 12.00 29.18 12.66 ;
    END
  END D[1]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 289.26 12.00 289.93 12.66 ;
      LAYER Metal6 ;
        RECT 289.26 12.00 289.93 12.66 ;
      LAYER Metal3 ;
        RECT 289.26 12.00 289.93 12.66 ;
      LAYER Metal4 ;
        RECT 289.26 12.00 289.93 12.66 ;
    END
  END D[20]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 297.31 12.00 297.96 12.66 ;
      LAYER Metal6 ;
        RECT 297.31 12.00 297.96 12.66 ;
      LAYER Metal3 ;
        RECT 297.31 12.00 297.96 12.66 ;
      LAYER Metal4 ;
        RECT 297.31 12.00 297.96 12.66 ;
    END
  END D[21]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 310.55 12.00 311.20 12.66 ;
      LAYER Metal6 ;
        RECT 310.55 12.00 311.20 12.66 ;
      LAYER Metal3 ;
        RECT 310.55 12.00 311.20 12.66 ;
      LAYER Metal4 ;
        RECT 310.55 12.00 311.20 12.66 ;
    END
  END D[22]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 318.58 12.00 319.25 12.66 ;
      LAYER Metal6 ;
        RECT 318.58 12.00 319.25 12.66 ;
      LAYER Metal3 ;
        RECT 318.58 12.00 319.25 12.66 ;
      LAYER Metal4 ;
        RECT 318.58 12.00 319.25 12.66 ;
    END
  END D[23]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 332.88 12.00 333.55 12.66 ;
      LAYER Metal6 ;
        RECT 332.88 12.00 333.55 12.66 ;
      LAYER Metal3 ;
        RECT 332.88 12.00 333.55 12.66 ;
      LAYER Metal4 ;
        RECT 332.88 12.00 333.55 12.66 ;
    END
  END D[24]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 340.93 12.00 341.58 12.66 ;
      LAYER Metal6 ;
        RECT 340.93 12.00 341.58 12.66 ;
      LAYER Metal3 ;
        RECT 340.93 12.00 341.58 12.66 ;
      LAYER Metal4 ;
        RECT 340.93 12.00 341.58 12.66 ;
    END
  END D[25]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 354.17 12.00 354.82 12.66 ;
      LAYER Metal6 ;
        RECT 354.17 12.00 354.82 12.66 ;
      LAYER Metal3 ;
        RECT 354.17 12.00 354.82 12.66 ;
      LAYER Metal4 ;
        RECT 354.17 12.00 354.82 12.66 ;
    END
  END D[26]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 362.20 12.00 362.87 12.66 ;
      LAYER Metal6 ;
        RECT 362.20 12.00 362.87 12.66 ;
      LAYER Metal3 ;
        RECT 362.20 12.00 362.87 12.66 ;
      LAYER Metal4 ;
        RECT 362.20 12.00 362.87 12.66 ;
    END
  END D[27]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.50 12.00 377.17 12.66 ;
      LAYER Metal6 ;
        RECT 376.50 12.00 377.17 12.66 ;
      LAYER Metal3 ;
        RECT 376.50 12.00 377.17 12.66 ;
      LAYER Metal4 ;
        RECT 376.50 12.00 377.17 12.66 ;
    END
  END D[28]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.55 12.00 385.20 12.66 ;
      LAYER Metal6 ;
        RECT 384.55 12.00 385.20 12.66 ;
      LAYER Metal3 ;
        RECT 384.55 12.00 385.20 12.66 ;
      LAYER Metal4 ;
        RECT 384.55 12.00 385.20 12.66 ;
    END
  END D[29]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 41.76 12.00 42.42 12.66 ;
      LAYER Metal6 ;
        RECT 41.76 12.00 42.42 12.66 ;
      LAYER Metal3 ;
        RECT 41.76 12.00 42.42 12.66 ;
      LAYER Metal4 ;
        RECT 41.76 12.00 42.42 12.66 ;
    END
  END D[2]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 397.79 12.00 398.44 12.66 ;
      LAYER Metal6 ;
        RECT 397.79 12.00 398.44 12.66 ;
      LAYER Metal3 ;
        RECT 397.79 12.00 398.44 12.66 ;
      LAYER Metal4 ;
        RECT 397.79 12.00 398.44 12.66 ;
    END
  END D[30]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 405.82 12.00 406.49 12.66 ;
      LAYER Metal6 ;
        RECT 405.82 12.00 406.49 12.66 ;
      LAYER Metal3 ;
        RECT 405.82 12.00 406.49 12.66 ;
      LAYER Metal4 ;
        RECT 405.82 12.00 406.49 12.66 ;
    END
  END D[31]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 49.80 12.00 50.46 12.66 ;
      LAYER Metal6 ;
        RECT 49.80 12.00 50.46 12.66 ;
      LAYER Metal3 ;
        RECT 49.80 12.00 50.46 12.66 ;
      LAYER Metal4 ;
        RECT 49.80 12.00 50.46 12.66 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.10 12.00 64.76 12.66 ;
      LAYER Metal6 ;
        RECT 64.10 12.00 64.76 12.66 ;
      LAYER Metal3 ;
        RECT 64.10 12.00 64.76 12.66 ;
      LAYER Metal4 ;
        RECT 64.10 12.00 64.76 12.66 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.14 12.00 72.80 12.66 ;
      LAYER Metal6 ;
        RECT 72.14 12.00 72.80 12.66 ;
      LAYER Metal3 ;
        RECT 72.14 12.00 72.80 12.66 ;
      LAYER Metal4 ;
        RECT 72.14 12.00 72.80 12.66 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.38 12.00 86.04 12.66 ;
      LAYER Metal6 ;
        RECT 85.38 12.00 86.04 12.66 ;
      LAYER Metal3 ;
        RECT 85.38 12.00 86.04 12.66 ;
      LAYER Metal4 ;
        RECT 85.38 12.00 86.04 12.66 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.42 12.00 94.08 12.66 ;
      LAYER Metal6 ;
        RECT 93.42 12.00 94.08 12.66 ;
      LAYER Metal3 ;
        RECT 93.42 12.00 94.08 12.66 ;
      LAYER Metal4 ;
        RECT 93.42 12.00 94.08 12.66 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.72 12.00 108.38 12.66 ;
      LAYER Metal6 ;
        RECT 107.72 12.00 108.38 12.66 ;
      LAYER Metal3 ;
        RECT 107.72 12.00 108.38 12.66 ;
      LAYER Metal4 ;
        RECT 107.72 12.00 108.38 12.66 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 115.76 12.00 116.42 12.66 ;
      LAYER Metal6 ;
        RECT 115.76 12.00 116.42 12.66 ;
      LAYER Metal3 ;
        RECT 115.76 12.00 116.42 12.66 ;
      LAYER Metal4 ;
        RECT 115.76 12.00 116.42 12.66 ;
    END
  END D[9]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 23.06 12.00 23.72 12.66 ;
      LAYER Metal6 ;
        RECT 23.06 12.00 23.72 12.66 ;
      LAYER Metal3 ;
        RECT 23.06 12.00 23.72 12.66 ;
      LAYER Metal4 ;
        RECT 23.06 12.00 23.72 12.66 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.58 12.00 132.24 12.66 ;
      LAYER Metal6 ;
        RECT 131.58 12.00 132.24 12.66 ;
      LAYER Metal3 ;
        RECT 131.58 12.00 132.24 12.66 ;
      LAYER Metal4 ;
        RECT 131.58 12.00 132.24 12.66 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 134.46 12.00 135.12 12.66 ;
      LAYER Metal6 ;
        RECT 134.46 12.00 135.12 12.66 ;
      LAYER Metal3 ;
        RECT 134.46 12.00 135.12 12.66 ;
      LAYER Metal4 ;
        RECT 134.46 12.00 135.12 12.66 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.92 12.00 154.58 12.66 ;
      LAYER Metal6 ;
        RECT 153.92 12.00 154.58 12.66 ;
      LAYER Metal3 ;
        RECT 153.92 12.00 154.58 12.66 ;
      LAYER Metal4 ;
        RECT 153.92 12.00 154.58 12.66 ;
    END
  END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 156.80 12.00 157.46 12.66 ;
      LAYER Metal6 ;
        RECT 156.80 12.00 157.46 12.66 ;
      LAYER Metal3 ;
        RECT 156.80 12.00 157.46 12.66 ;
      LAYER Metal4 ;
        RECT 156.80 12.00 157.46 12.66 ;
    END
  END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.20 12.00 175.86 12.66 ;
      LAYER Metal6 ;
        RECT 175.20 12.00 175.86 12.66 ;
      LAYER Metal3 ;
        RECT 175.20 12.00 175.86 12.66 ;
      LAYER Metal4 ;
        RECT 175.20 12.00 175.86 12.66 ;
    END
  END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.08 12.00 178.74 12.66 ;
      LAYER Metal6 ;
        RECT 178.08 12.00 178.74 12.66 ;
      LAYER Metal3 ;
        RECT 178.08 12.00 178.74 12.66 ;
      LAYER Metal4 ;
        RECT 178.08 12.00 178.74 12.66 ;
    END
  END Q[15]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 248.22 12.00 248.88 12.66 ;
      LAYER Metal6 ;
        RECT 248.22 12.00 248.88 12.66 ;
      LAYER Metal3 ;
        RECT 248.22 12.00 248.88 12.66 ;
      LAYER Metal4 ;
        RECT 248.22 12.00 248.88 12.66 ;
    END
  END Q[16]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 251.10 12.00 251.76 12.66 ;
      LAYER Metal6 ;
        RECT 251.10 12.00 251.76 12.66 ;
      LAYER Metal3 ;
        RECT 251.10 12.00 251.76 12.66 ;
      LAYER Metal4 ;
        RECT 251.10 12.00 251.76 12.66 ;
    END
  END Q[17]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 269.50 12.00 270.17 12.66 ;
      LAYER Metal6 ;
        RECT 269.50 12.00 270.17 12.66 ;
      LAYER Metal3 ;
        RECT 269.50 12.00 270.17 12.66 ;
      LAYER Metal4 ;
        RECT 269.50 12.00 270.17 12.66 ;
    END
  END Q[18]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 272.38 12.00 273.05 12.66 ;
      LAYER Metal6 ;
        RECT 272.38 12.00 273.05 12.66 ;
      LAYER Metal3 ;
        RECT 272.38 12.00 273.05 12.66 ;
      LAYER Metal4 ;
        RECT 272.38 12.00 273.05 12.66 ;
    END
  END Q[19]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.94 12.00 26.60 12.66 ;
      LAYER Metal6 ;
        RECT 25.94 12.00 26.60 12.66 ;
      LAYER Metal3 ;
        RECT 25.94 12.00 26.60 12.66 ;
      LAYER Metal4 ;
        RECT 25.94 12.00 26.60 12.66 ;
    END
  END Q[1]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.85 12.00 292.50 12.66 ;
      LAYER Metal6 ;
        RECT 291.85 12.00 292.50 12.66 ;
      LAYER Metal3 ;
        RECT 291.85 12.00 292.50 12.66 ;
      LAYER Metal4 ;
        RECT 291.85 12.00 292.50 12.66 ;
    END
  END Q[20]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 294.73 12.00 295.38 12.66 ;
      LAYER Metal6 ;
        RECT 294.73 12.00 295.38 12.66 ;
      LAYER Metal3 ;
        RECT 294.73 12.00 295.38 12.66 ;
      LAYER Metal4 ;
        RECT 294.73 12.00 295.38 12.66 ;
    END
  END Q[21]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 313.12 12.00 313.79 12.66 ;
      LAYER Metal6 ;
        RECT 313.12 12.00 313.79 12.66 ;
      LAYER Metal3 ;
        RECT 313.12 12.00 313.79 12.66 ;
      LAYER Metal4 ;
        RECT 313.12 12.00 313.79 12.66 ;
    END
  END Q[22]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 316.00 12.00 316.67 12.66 ;
      LAYER Metal6 ;
        RECT 316.00 12.00 316.67 12.66 ;
      LAYER Metal3 ;
        RECT 316.00 12.00 316.67 12.66 ;
      LAYER Metal4 ;
        RECT 316.00 12.00 316.67 12.66 ;
    END
  END Q[23]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 335.46 12.00 336.12 12.66 ;
      LAYER Metal6 ;
        RECT 335.46 12.00 336.12 12.66 ;
      LAYER Metal3 ;
        RECT 335.46 12.00 336.12 12.66 ;
      LAYER Metal4 ;
        RECT 335.46 12.00 336.12 12.66 ;
    END
  END Q[24]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 338.35 12.00 339.00 12.66 ;
      LAYER Metal6 ;
        RECT 338.35 12.00 339.00 12.66 ;
      LAYER Metal3 ;
        RECT 338.35 12.00 339.00 12.66 ;
      LAYER Metal4 ;
        RECT 338.35 12.00 339.00 12.66 ;
    END
  END Q[25]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 356.75 12.00 357.40 12.66 ;
      LAYER Metal6 ;
        RECT 356.75 12.00 357.40 12.66 ;
      LAYER Metal3 ;
        RECT 356.75 12.00 357.40 12.66 ;
      LAYER Metal4 ;
        RECT 356.75 12.00 357.40 12.66 ;
    END
  END Q[26]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 359.62 12.00 360.29 12.66 ;
      LAYER Metal6 ;
        RECT 359.62 12.00 360.29 12.66 ;
      LAYER Metal3 ;
        RECT 359.62 12.00 360.29 12.66 ;
      LAYER Metal4 ;
        RECT 359.62 12.00 360.29 12.66 ;
    END
  END Q[27]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 379.08 12.00 379.75 12.66 ;
      LAYER Metal6 ;
        RECT 379.08 12.00 379.75 12.66 ;
      LAYER Metal3 ;
        RECT 379.08 12.00 379.75 12.66 ;
      LAYER Metal4 ;
        RECT 379.08 12.00 379.75 12.66 ;
    END
  END Q[28]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 381.96 12.00 382.62 12.66 ;
      LAYER Metal6 ;
        RECT 381.96 12.00 382.62 12.66 ;
      LAYER Metal3 ;
        RECT 381.96 12.00 382.62 12.66 ;
      LAYER Metal4 ;
        RECT 381.96 12.00 382.62 12.66 ;
    END
  END Q[29]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 44.34 12.00 45.00 12.66 ;
      LAYER Metal6 ;
        RECT 44.34 12.00 45.00 12.66 ;
      LAYER Metal3 ;
        RECT 44.34 12.00 45.00 12.66 ;
      LAYER Metal4 ;
        RECT 44.34 12.00 45.00 12.66 ;
    END
  END Q[2]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 400.37 12.00 401.02 12.66 ;
      LAYER Metal6 ;
        RECT 400.37 12.00 401.02 12.66 ;
      LAYER Metal3 ;
        RECT 400.37 12.00 401.02 12.66 ;
      LAYER Metal4 ;
        RECT 400.37 12.00 401.02 12.66 ;
    END
  END Q[30]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 403.25 12.00 403.90 12.66 ;
      LAYER Metal6 ;
        RECT 403.25 12.00 403.90 12.66 ;
      LAYER Metal3 ;
        RECT 403.25 12.00 403.90 12.66 ;
      LAYER Metal4 ;
        RECT 403.25 12.00 403.90 12.66 ;
    END
  END Q[31]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.22 12.00 47.88 12.66 ;
      LAYER Metal6 ;
        RECT 47.22 12.00 47.88 12.66 ;
      LAYER Metal3 ;
        RECT 47.22 12.00 47.88 12.66 ;
      LAYER Metal4 ;
        RECT 47.22 12.00 47.88 12.66 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 66.68 12.00 67.34 12.66 ;
      LAYER Metal6 ;
        RECT 66.68 12.00 67.34 12.66 ;
      LAYER Metal3 ;
        RECT 66.68 12.00 67.34 12.66 ;
      LAYER Metal4 ;
        RECT 66.68 12.00 67.34 12.66 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.56 12.00 70.22 12.66 ;
      LAYER Metal6 ;
        RECT 69.56 12.00 70.22 12.66 ;
      LAYER Metal3 ;
        RECT 69.56 12.00 70.22 12.66 ;
      LAYER Metal4 ;
        RECT 69.56 12.00 70.22 12.66 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 87.96 12.00 88.62 12.66 ;
      LAYER Metal6 ;
        RECT 87.96 12.00 88.62 12.66 ;
      LAYER Metal3 ;
        RECT 87.96 12.00 88.62 12.66 ;
      LAYER Metal4 ;
        RECT 87.96 12.00 88.62 12.66 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.84 12.00 91.50 12.66 ;
      LAYER Metal6 ;
        RECT 90.84 12.00 91.50 12.66 ;
      LAYER Metal3 ;
        RECT 90.84 12.00 91.50 12.66 ;
      LAYER Metal4 ;
        RECT 90.84 12.00 91.50 12.66 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.30 12.00 110.96 12.66 ;
      LAYER Metal6 ;
        RECT 110.30 12.00 110.96 12.66 ;
      LAYER Metal3 ;
        RECT 110.30 12.00 110.96 12.66 ;
      LAYER Metal4 ;
        RECT 110.30 12.00 110.96 12.66 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 113.18 12.00 113.84 12.66 ;
      LAYER Metal6 ;
        RECT 113.18 12.00 113.84 12.66 ;
      LAYER Metal3 ;
        RECT 113.18 12.00 113.84 12.66 ;
      LAYER Metal4 ;
        RECT 113.18 12.00 113.84 12.66 ;
    END
  END Q[9]
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 234.48 12.00 235.14 12.66 ;
      LAYER Metal6 ;
        RECT 234.48 12.00 235.14 12.66 ;
      LAYER Metal3 ;
        RECT 234.48 12.00 235.14 12.66 ;
      LAYER Metal4 ;
        RECT 234.48 12.00 235.14 12.66 ;
    END
  END WE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 109.22 426.96 114.22 ;
        RECT 0.00 0.00 426.96 5.00 ;
      LAYER Metal2 ;
        RECT 421.96 0.00 426.96 114.22 ;
        RECT 0.00 0.00 5.00 114.22 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.60 103.61 421.37 108.61 ;
        RECT 5.60 5.60 421.37 10.60 ;
      LAYER Metal2 ;
        RECT 416.37 5.60 421.37 108.61 ;
        RECT 5.60 5.60 10.60 108.61 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12.00 12.00 415.01 102.02 ;
    LAYER Metal2 ;
      RECT 12.00 12.00 415.01 102.02 ;
    LAYER Metal3 ;
      RECT 12.00 12.00 415.01 102.02 ;
    LAYER Metal4 ;
      RECT 12.00 12.00 415.01 102.02 ;
    LAYER Metal5 ;
      RECT 12.00 12.00 415.01 102.02 ;
    LAYER Metal6 ;
      RECT 12.00 12.00 415.01 102.02 ;
  END
END MEM1

MACRO MEM2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2 0 0 ;
  SIZE 423.015 BY 145.035 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 102.42 12.66 103.08 ;
      LAYER Metal6 ;
        RECT 12.00 102.42 12.66 103.08 ;
      LAYER Metal3 ;
        RECT 12.00 102.42 12.66 103.08 ;
      LAYER Metal4 ;
        RECT 12.00 102.42 12.66 103.08 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 96.30 12.66 96.96 ;
      LAYER Metal6 ;
        RECT 12.00 96.30 12.66 96.96 ;
      LAYER Metal3 ;
        RECT 12.00 96.30 12.66 96.96 ;
      LAYER Metal4 ;
        RECT 12.00 96.30 12.66 96.96 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 87.08 12.66 87.74 ;
      LAYER Metal6 ;
        RECT 12.00 87.08 12.66 87.74 ;
      LAYER Metal3 ;
        RECT 12.00 87.08 12.66 87.74 ;
      LAYER Metal4 ;
        RECT 12.00 87.08 12.66 87.74 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 84.06 12.66 84.72 ;
      LAYER Metal6 ;
        RECT 12.00 84.06 12.66 84.72 ;
      LAYER Metal3 ;
        RECT 12.00 84.06 12.66 84.72 ;
      LAYER Metal4 ;
        RECT 12.00 84.06 12.66 84.72 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 80.96 12.66 81.62 ;
      LAYER Metal6 ;
        RECT 12.00 80.96 12.66 81.62 ;
      LAYER Metal3 ;
        RECT 12.00 80.96 12.66 81.62 ;
      LAYER Metal4 ;
        RECT 12.00 80.96 12.66 81.62 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 74.84 12.66 75.50 ;
      LAYER Metal6 ;
        RECT 12.00 74.84 12.66 75.50 ;
      LAYER Metal3 ;
        RECT 12.00 74.84 12.66 75.50 ;
      LAYER Metal4 ;
        RECT 12.00 74.84 12.66 75.50 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 71.82 12.66 72.48 ;
      LAYER Metal6 ;
        RECT 12.00 71.82 12.66 72.48 ;
      LAYER Metal3 ;
        RECT 12.00 71.82 12.66 72.48 ;
      LAYER Metal4 ;
        RECT 12.00 71.82 12.66 72.48 ;
    END
  END A1[6]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 36.40 12.66 37.06 ;
      LAYER Metal6 ;
        RECT 12.00 36.40 12.66 37.06 ;
      LAYER Metal3 ;
        RECT 12.00 36.40 12.66 37.06 ;
      LAYER Metal4 ;
        RECT 12.00 36.40 12.66 37.06 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 42.52 12.66 43.18 ;
      LAYER Metal6 ;
        RECT 12.00 42.52 12.66 43.18 ;
      LAYER Metal3 ;
        RECT 12.00 42.52 12.66 43.18 ;
      LAYER Metal4 ;
        RECT 12.00 42.52 12.66 43.18 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 51.74 12.66 52.40 ;
      LAYER Metal6 ;
        RECT 12.00 51.74 12.66 52.40 ;
      LAYER Metal3 ;
        RECT 12.00 51.74 12.66 52.40 ;
      LAYER Metal4 ;
        RECT 12.00 51.74 12.66 52.40 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 54.76 12.66 55.42 ;
      LAYER Metal6 ;
        RECT 12.00 54.76 12.66 55.42 ;
      LAYER Metal3 ;
        RECT 12.00 54.76 12.66 55.42 ;
      LAYER Metal4 ;
        RECT 12.00 54.76 12.66 55.42 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 57.86 12.66 58.52 ;
      LAYER Metal6 ;
        RECT 12.00 57.86 12.66 58.52 ;
      LAYER Metal3 ;
        RECT 12.00 57.86 12.66 58.52 ;
      LAYER Metal4 ;
        RECT 12.00 57.86 12.66 58.52 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 63.98 12.66 64.64 ;
      LAYER Metal6 ;
        RECT 12.00 63.98 12.66 64.64 ;
      LAYER Metal3 ;
        RECT 12.00 63.98 12.66 64.64 ;
      LAYER Metal4 ;
        RECT 12.00 63.98 12.66 64.64 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 67.00 12.66 67.66 ;
      LAYER Metal6 ;
        RECT 12.00 67.00 12.66 67.66 ;
      LAYER Metal3 ;
        RECT 12.00 67.00 12.66 67.66 ;
      LAYER Metal4 ;
        RECT 12.00 67.00 12.66 67.66 ;
    END
  END A2[6]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 210.28 12.00 210.94 12.66 ;
      LAYER Metal6 ;
        RECT 210.28 12.00 210.94 12.66 ;
      LAYER Metal3 ;
        RECT 210.28 12.00 210.94 12.66 ;
      LAYER Metal4 ;
        RECT 210.28 12.00 210.94 12.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 196.36 12.00 197.02 12.66 ;
      LAYER Metal6 ;
        RECT 196.36 12.00 197.02 12.66 ;
      LAYER Metal3 ;
        RECT 196.36 12.00 197.02 12.66 ;
      LAYER Metal4 ;
        RECT 196.36 12.00 197.02 12.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 218.91 12.00 219.56 12.66 ;
      LAYER Metal6 ;
        RECT 218.91 12.00 219.56 12.66 ;
      LAYER Metal3 ;
        RECT 218.91 12.00 219.56 12.66 ;
      LAYER Metal4 ;
        RECT 218.91 12.00 219.56 12.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 187.74 12.00 188.40 12.66 ;
      LAYER Metal6 ;
        RECT 187.74 12.00 188.40 12.66 ;
      LAYER Metal3 ;
        RECT 187.74 12.00 188.40 12.66 ;
      LAYER Metal4 ;
        RECT 187.74 12.00 188.40 12.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 15.86 12.00 16.52 12.66 ;
      LAYER Metal6 ;
        RECT 15.86 12.00 16.52 12.66 ;
      LAYER Metal3 ;
        RECT 15.86 12.00 16.52 12.66 ;
      LAYER Metal4 ;
        RECT 15.86 12.00 16.52 12.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 122.26 12.00 122.92 12.66 ;
      LAYER Metal6 ;
        RECT 122.26 12.00 122.92 12.66 ;
      LAYER Metal3 ;
        RECT 122.26 12.00 122.92 12.66 ;
      LAYER Metal4 ;
        RECT 122.26 12.00 122.92 12.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 142.40 12.00 143.06 12.66 ;
      LAYER Metal6 ;
        RECT 142.40 12.00 143.06 12.66 ;
      LAYER Metal3 ;
        RECT 142.40 12.00 143.06 12.66 ;
      LAYER Metal4 ;
        RECT 142.40 12.00 143.06 12.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 143.54 12.00 144.20 12.66 ;
      LAYER Metal6 ;
        RECT 143.54 12.00 144.20 12.66 ;
      LAYER Metal3 ;
        RECT 143.54 12.00 144.20 12.66 ;
      LAYER Metal4 ;
        RECT 143.54 12.00 144.20 12.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 163.68 12.00 164.34 12.66 ;
      LAYER Metal6 ;
        RECT 163.68 12.00 164.34 12.66 ;
      LAYER Metal3 ;
        RECT 163.68 12.00 164.34 12.66 ;
      LAYER Metal4 ;
        RECT 163.68 12.00 164.34 12.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 164.82 12.00 165.48 12.66 ;
      LAYER Metal6 ;
        RECT 164.82 12.00 165.48 12.66 ;
      LAYER Metal3 ;
        RECT 164.82 12.00 165.48 12.66 ;
      LAYER Metal4 ;
        RECT 164.82 12.00 165.48 12.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 184.96 12.00 185.62 12.66 ;
      LAYER Metal6 ;
        RECT 184.96 12.00 185.62 12.66 ;
      LAYER Metal3 ;
        RECT 184.96 12.00 185.62 12.66 ;
      LAYER Metal4 ;
        RECT 184.96 12.00 185.62 12.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 221.68 12.00 222.34 12.66 ;
      LAYER Metal6 ;
        RECT 221.68 12.00 222.34 12.66 ;
      LAYER Metal3 ;
        RECT 221.68 12.00 222.34 12.66 ;
      LAYER Metal4 ;
        RECT 221.68 12.00 222.34 12.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 241.82 12.00 242.48 12.66 ;
      LAYER Metal6 ;
        RECT 241.82 12.00 242.48 12.66 ;
      LAYER Metal3 ;
        RECT 241.82 12.00 242.48 12.66 ;
      LAYER Metal4 ;
        RECT 241.82 12.00 242.48 12.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 242.96 12.00 243.62 12.66 ;
      LAYER Metal6 ;
        RECT 242.96 12.00 243.62 12.66 ;
      LAYER Metal3 ;
        RECT 242.96 12.00 243.62 12.66 ;
      LAYER Metal4 ;
        RECT 242.96 12.00 243.62 12.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 263.10 12.00 263.76 12.66 ;
      LAYER Metal6 ;
        RECT 263.10 12.00 263.76 12.66 ;
      LAYER Metal3 ;
        RECT 263.10 12.00 263.76 12.66 ;
      LAYER Metal4 ;
        RECT 263.10 12.00 263.76 12.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 36.00 12.00 36.66 12.66 ;
      LAYER Metal6 ;
        RECT 36.00 12.00 36.66 12.66 ;
      LAYER Metal3 ;
        RECT 36.00 12.00 36.66 12.66 ;
      LAYER Metal4 ;
        RECT 36.00 12.00 36.66 12.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 264.24 12.00 264.90 12.66 ;
      LAYER Metal6 ;
        RECT 264.24 12.00 264.90 12.66 ;
      LAYER Metal3 ;
        RECT 264.24 12.00 264.90 12.66 ;
      LAYER Metal4 ;
        RECT 264.24 12.00 264.90 12.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 284.38 12.00 285.04 12.66 ;
      LAYER Metal6 ;
        RECT 284.38 12.00 285.04 12.66 ;
      LAYER Metal3 ;
        RECT 284.38 12.00 285.04 12.66 ;
      LAYER Metal4 ;
        RECT 284.38 12.00 285.04 12.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 285.52 12.00 286.18 12.66 ;
      LAYER Metal6 ;
        RECT 285.52 12.00 286.18 12.66 ;
      LAYER Metal3 ;
        RECT 285.52 12.00 286.18 12.66 ;
      LAYER Metal4 ;
        RECT 285.52 12.00 286.18 12.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 305.66 12.00 306.32 12.66 ;
      LAYER Metal6 ;
        RECT 305.66 12.00 306.32 12.66 ;
      LAYER Metal3 ;
        RECT 305.66 12.00 306.32 12.66 ;
      LAYER Metal4 ;
        RECT 305.66 12.00 306.32 12.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 306.80 12.00 307.46 12.66 ;
      LAYER Metal6 ;
        RECT 306.80 12.00 307.46 12.66 ;
      LAYER Metal3 ;
        RECT 306.80 12.00 307.46 12.66 ;
      LAYER Metal4 ;
        RECT 306.80 12.00 307.46 12.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 326.94 12.00 327.60 12.66 ;
      LAYER Metal6 ;
        RECT 326.94 12.00 327.60 12.66 ;
      LAYER Metal3 ;
        RECT 326.94 12.00 327.60 12.66 ;
      LAYER Metal4 ;
        RECT 326.94 12.00 327.60 12.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 328.08 12.00 328.74 12.66 ;
      LAYER Metal6 ;
        RECT 328.08 12.00 328.74 12.66 ;
      LAYER Metal3 ;
        RECT 328.08 12.00 328.74 12.66 ;
      LAYER Metal4 ;
        RECT 328.08 12.00 328.74 12.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 348.22 12.00 348.88 12.66 ;
      LAYER Metal6 ;
        RECT 348.22 12.00 348.88 12.66 ;
      LAYER Metal3 ;
        RECT 348.22 12.00 348.88 12.66 ;
      LAYER Metal4 ;
        RECT 348.22 12.00 348.88 12.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 349.36 12.00 350.02 12.66 ;
      LAYER Metal6 ;
        RECT 349.36 12.00 350.02 12.66 ;
      LAYER Metal3 ;
        RECT 349.36 12.00 350.02 12.66 ;
      LAYER Metal4 ;
        RECT 349.36 12.00 350.02 12.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 369.50 12.00 370.16 12.66 ;
      LAYER Metal6 ;
        RECT 369.50 12.00 370.16 12.66 ;
      LAYER Metal3 ;
        RECT 369.50 12.00 370.16 12.66 ;
      LAYER Metal4 ;
        RECT 369.50 12.00 370.16 12.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 37.14 12.00 37.80 12.66 ;
      LAYER Metal6 ;
        RECT 37.14 12.00 37.80 12.66 ;
      LAYER Metal3 ;
        RECT 37.14 12.00 37.80 12.66 ;
      LAYER Metal4 ;
        RECT 37.14 12.00 37.80 12.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 370.64 12.00 371.30 12.66 ;
      LAYER Metal6 ;
        RECT 370.64 12.00 371.30 12.66 ;
      LAYER Metal3 ;
        RECT 370.64 12.00 371.30 12.66 ;
      LAYER Metal4 ;
        RECT 370.64 12.00 371.30 12.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 390.78 12.00 391.44 12.66 ;
      LAYER Metal6 ;
        RECT 390.78 12.00 391.44 12.66 ;
      LAYER Metal3 ;
        RECT 390.78 12.00 391.44 12.66 ;
      LAYER Metal4 ;
        RECT 390.78 12.00 391.44 12.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 57.28 12.00 57.94 12.66 ;
      LAYER Metal6 ;
        RECT 57.28 12.00 57.94 12.66 ;
      LAYER Metal3 ;
        RECT 57.28 12.00 57.94 12.66 ;
      LAYER Metal4 ;
        RECT 57.28 12.00 57.94 12.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 58.42 12.00 59.08 12.66 ;
      LAYER Metal6 ;
        RECT 58.42 12.00 59.08 12.66 ;
      LAYER Metal3 ;
        RECT 58.42 12.00 59.08 12.66 ;
      LAYER Metal4 ;
        RECT 58.42 12.00 59.08 12.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 78.56 12.00 79.22 12.66 ;
      LAYER Metal6 ;
        RECT 78.56 12.00 79.22 12.66 ;
      LAYER Metal3 ;
        RECT 78.56 12.00 79.22 12.66 ;
      LAYER Metal4 ;
        RECT 78.56 12.00 79.22 12.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 79.70 12.00 80.36 12.66 ;
      LAYER Metal6 ;
        RECT 79.70 12.00 80.36 12.66 ;
      LAYER Metal3 ;
        RECT 79.70 12.00 80.36 12.66 ;
      LAYER Metal4 ;
        RECT 79.70 12.00 80.36 12.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 99.84 12.00 100.50 12.66 ;
      LAYER Metal6 ;
        RECT 99.84 12.00 100.50 12.66 ;
      LAYER Metal3 ;
        RECT 99.84 12.00 100.50 12.66 ;
      LAYER Metal4 ;
        RECT 99.84 12.00 100.50 12.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 100.98 12.00 101.64 12.66 ;
      LAYER Metal6 ;
        RECT 100.98 12.00 101.64 12.66 ;
      LAYER Metal3 ;
        RECT 100.98 12.00 101.64 12.66 ;
      LAYER Metal4 ;
        RECT 100.98 12.00 101.64 12.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 121.12 12.00 121.78 12.66 ;
      LAYER Metal6 ;
        RECT 121.12 12.00 121.78 12.66 ;
      LAYER Metal3 ;
        RECT 121.12 12.00 121.78 12.66 ;
      LAYER Metal4 ;
        RECT 121.12 12.00 121.78 12.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.36 12.00 26.02 12.66 ;
      LAYER Metal6 ;
        RECT 25.36 12.00 26.02 12.66 ;
      LAYER Metal3 ;
        RECT 25.36 12.00 26.02 12.66 ;
      LAYER Metal4 ;
        RECT 25.36 12.00 26.02 12.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.76 12.00 132.42 12.66 ;
      LAYER Metal6 ;
        RECT 131.76 12.00 132.42 12.66 ;
      LAYER Metal3 ;
        RECT 131.76 12.00 132.42 12.66 ;
      LAYER Metal4 ;
        RECT 131.76 12.00 132.42 12.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 132.90 12.00 133.56 12.66 ;
      LAYER Metal6 ;
        RECT 132.90 12.00 133.56 12.66 ;
      LAYER Metal3 ;
        RECT 132.90 12.00 133.56 12.66 ;
      LAYER Metal4 ;
        RECT 132.90 12.00 133.56 12.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.04 12.00 153.70 12.66 ;
      LAYER Metal6 ;
        RECT 153.04 12.00 153.70 12.66 ;
      LAYER Metal3 ;
        RECT 153.04 12.00 153.70 12.66 ;
      LAYER Metal4 ;
        RECT 153.04 12.00 153.70 12.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 154.18 12.00 154.84 12.66 ;
      LAYER Metal6 ;
        RECT 154.18 12.00 154.84 12.66 ;
      LAYER Metal3 ;
        RECT 154.18 12.00 154.84 12.66 ;
      LAYER Metal4 ;
        RECT 154.18 12.00 154.84 12.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 174.32 12.00 174.98 12.66 ;
      LAYER Metal6 ;
        RECT 174.32 12.00 174.98 12.66 ;
      LAYER Metal3 ;
        RECT 174.32 12.00 174.98 12.66 ;
      LAYER Metal4 ;
        RECT 174.32 12.00 174.98 12.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.46 12.00 176.12 12.66 ;
      LAYER Metal6 ;
        RECT 175.46 12.00 176.12 12.66 ;
      LAYER Metal3 ;
        RECT 175.46 12.00 176.12 12.66 ;
      LAYER Metal4 ;
        RECT 175.46 12.00 176.12 12.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 231.18 12.00 231.84 12.66 ;
      LAYER Metal6 ;
        RECT 231.18 12.00 231.84 12.66 ;
      LAYER Metal3 ;
        RECT 231.18 12.00 231.84 12.66 ;
      LAYER Metal4 ;
        RECT 231.18 12.00 231.84 12.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 232.32 12.00 232.98 12.66 ;
      LAYER Metal6 ;
        RECT 232.32 12.00 232.98 12.66 ;
      LAYER Metal3 ;
        RECT 232.32 12.00 232.98 12.66 ;
      LAYER Metal4 ;
        RECT 232.32 12.00 232.98 12.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 252.46 12.00 253.12 12.66 ;
      LAYER Metal6 ;
        RECT 252.46 12.00 253.12 12.66 ;
      LAYER Metal3 ;
        RECT 252.46 12.00 253.12 12.66 ;
      LAYER Metal4 ;
        RECT 252.46 12.00 253.12 12.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 253.60 12.00 254.26 12.66 ;
      LAYER Metal6 ;
        RECT 253.60 12.00 254.26 12.66 ;
      LAYER Metal3 ;
        RECT 253.60 12.00 254.26 12.66 ;
      LAYER Metal4 ;
        RECT 253.60 12.00 254.26 12.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 26.50 12.00 27.16 12.66 ;
      LAYER Metal6 ;
        RECT 26.50 12.00 27.16 12.66 ;
      LAYER Metal3 ;
        RECT 26.50 12.00 27.16 12.66 ;
      LAYER Metal4 ;
        RECT 26.50 12.00 27.16 12.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 273.74 12.00 274.40 12.66 ;
      LAYER Metal6 ;
        RECT 273.74 12.00 274.40 12.66 ;
      LAYER Metal3 ;
        RECT 273.74 12.00 274.40 12.66 ;
      LAYER Metal4 ;
        RECT 273.74 12.00 274.40 12.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 274.88 12.00 275.54 12.66 ;
      LAYER Metal6 ;
        RECT 274.88 12.00 275.54 12.66 ;
      LAYER Metal3 ;
        RECT 274.88 12.00 275.54 12.66 ;
      LAYER Metal4 ;
        RECT 274.88 12.00 275.54 12.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 295.02 12.00 295.68 12.66 ;
      LAYER Metal6 ;
        RECT 295.02 12.00 295.68 12.66 ;
      LAYER Metal3 ;
        RECT 295.02 12.00 295.68 12.66 ;
      LAYER Metal4 ;
        RECT 295.02 12.00 295.68 12.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 296.16 12.00 296.82 12.66 ;
      LAYER Metal6 ;
        RECT 296.16 12.00 296.82 12.66 ;
      LAYER Metal3 ;
        RECT 296.16 12.00 296.82 12.66 ;
      LAYER Metal4 ;
        RECT 296.16 12.00 296.82 12.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 316.30 12.00 316.96 12.66 ;
      LAYER Metal6 ;
        RECT 316.30 12.00 316.96 12.66 ;
      LAYER Metal3 ;
        RECT 316.30 12.00 316.96 12.66 ;
      LAYER Metal4 ;
        RECT 316.30 12.00 316.96 12.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 317.44 12.00 318.10 12.66 ;
      LAYER Metal6 ;
        RECT 317.44 12.00 318.10 12.66 ;
      LAYER Metal3 ;
        RECT 317.44 12.00 318.10 12.66 ;
      LAYER Metal4 ;
        RECT 317.44 12.00 318.10 12.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 337.58 12.00 338.24 12.66 ;
      LAYER Metal6 ;
        RECT 337.58 12.00 338.24 12.66 ;
      LAYER Metal3 ;
        RECT 337.58 12.00 338.24 12.66 ;
      LAYER Metal4 ;
        RECT 337.58 12.00 338.24 12.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 338.72 12.00 339.38 12.66 ;
      LAYER Metal6 ;
        RECT 338.72 12.00 339.38 12.66 ;
      LAYER Metal3 ;
        RECT 338.72 12.00 339.38 12.66 ;
      LAYER Metal4 ;
        RECT 338.72 12.00 339.38 12.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 358.86 12.00 359.52 12.66 ;
      LAYER Metal6 ;
        RECT 358.86 12.00 359.52 12.66 ;
      LAYER Metal3 ;
        RECT 358.86 12.00 359.52 12.66 ;
      LAYER Metal4 ;
        RECT 358.86 12.00 359.52 12.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 360.00 12.00 360.66 12.66 ;
      LAYER Metal6 ;
        RECT 360.00 12.00 360.66 12.66 ;
      LAYER Metal3 ;
        RECT 360.00 12.00 360.66 12.66 ;
      LAYER Metal4 ;
        RECT 360.00 12.00 360.66 12.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 46.64 12.00 47.30 12.66 ;
      LAYER Metal6 ;
        RECT 46.64 12.00 47.30 12.66 ;
      LAYER Metal3 ;
        RECT 46.64 12.00 47.30 12.66 ;
      LAYER Metal4 ;
        RECT 46.64 12.00 47.30 12.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 380.14 12.00 380.80 12.66 ;
      LAYER Metal6 ;
        RECT 380.14 12.00 380.80 12.66 ;
      LAYER Metal3 ;
        RECT 380.14 12.00 380.80 12.66 ;
      LAYER Metal4 ;
        RECT 380.14 12.00 380.80 12.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 381.28 12.00 381.94 12.66 ;
      LAYER Metal6 ;
        RECT 381.28 12.00 381.94 12.66 ;
      LAYER Metal3 ;
        RECT 381.28 12.00 381.94 12.66 ;
      LAYER Metal4 ;
        RECT 381.28 12.00 381.94 12.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.78 12.00 48.44 12.66 ;
      LAYER Metal6 ;
        RECT 47.78 12.00 48.44 12.66 ;
      LAYER Metal3 ;
        RECT 47.78 12.00 48.44 12.66 ;
      LAYER Metal4 ;
        RECT 47.78 12.00 48.44 12.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 67.92 12.00 68.58 12.66 ;
      LAYER Metal6 ;
        RECT 67.92 12.00 68.58 12.66 ;
      LAYER Metal3 ;
        RECT 67.92 12.00 68.58 12.66 ;
      LAYER Metal4 ;
        RECT 67.92 12.00 68.58 12.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.06 12.00 69.72 12.66 ;
      LAYER Metal6 ;
        RECT 69.06 12.00 69.72 12.66 ;
      LAYER Metal3 ;
        RECT 69.06 12.00 69.72 12.66 ;
      LAYER Metal4 ;
        RECT 69.06 12.00 69.72 12.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 89.20 12.00 89.86 12.66 ;
      LAYER Metal6 ;
        RECT 89.20 12.00 89.86 12.66 ;
      LAYER Metal3 ;
        RECT 89.20 12.00 89.86 12.66 ;
      LAYER Metal4 ;
        RECT 89.20 12.00 89.86 12.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.34 12.00 91.00 12.66 ;
      LAYER Metal6 ;
        RECT 90.34 12.00 91.00 12.66 ;
      LAYER Metal3 ;
        RECT 90.34 12.00 91.00 12.66 ;
      LAYER Metal4 ;
        RECT 90.34 12.00 91.00 12.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.48 12.00 111.14 12.66 ;
      LAYER Metal6 ;
        RECT 110.48 12.00 111.14 12.66 ;
      LAYER Metal3 ;
        RECT 110.48 12.00 111.14 12.66 ;
      LAYER Metal4 ;
        RECT 110.48 12.00 111.14 12.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 111.62 12.00 112.28 12.66 ;
      LAYER Metal6 ;
        RECT 111.62 12.00 112.28 12.66 ;
      LAYER Metal3 ;
        RECT 111.62 12.00 112.28 12.66 ;
      LAYER Metal4 ;
        RECT 111.62 12.00 112.28 12.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 18.28 12.00 18.94 12.66 ;
      LAYER Metal6 ;
        RECT 18.28 12.00 18.94 12.66 ;
      LAYER Metal3 ;
        RECT 18.28 12.00 18.94 12.66 ;
      LAYER Metal4 ;
        RECT 18.28 12.00 18.94 12.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 125.56 12.00 126.22 12.66 ;
      LAYER Metal6 ;
        RECT 125.56 12.00 126.22 12.66 ;
      LAYER Metal3 ;
        RECT 125.56 12.00 126.22 12.66 ;
      LAYER Metal4 ;
        RECT 125.56 12.00 126.22 12.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 139.10 12.00 139.76 12.66 ;
      LAYER Metal6 ;
        RECT 139.10 12.00 139.76 12.66 ;
      LAYER Metal3 ;
        RECT 139.10 12.00 139.76 12.66 ;
      LAYER Metal4 ;
        RECT 139.10 12.00 139.76 12.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 146.84 12.00 147.50 12.66 ;
      LAYER Metal6 ;
        RECT 146.84 12.00 147.50 12.66 ;
      LAYER Metal3 ;
        RECT 146.84 12.00 147.50 12.66 ;
      LAYER Metal4 ;
        RECT 146.84 12.00 147.50 12.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 160.38 12.00 161.04 12.66 ;
      LAYER Metal6 ;
        RECT 160.38 12.00 161.04 12.66 ;
      LAYER Metal3 ;
        RECT 160.38 12.00 161.04 12.66 ;
      LAYER Metal4 ;
        RECT 160.38 12.00 161.04 12.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 168.12 12.00 168.78 12.66 ;
      LAYER Metal6 ;
        RECT 168.12 12.00 168.78 12.66 ;
      LAYER Metal3 ;
        RECT 168.12 12.00 168.78 12.66 ;
      LAYER Metal4 ;
        RECT 168.12 12.00 168.78 12.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 181.66 12.00 182.32 12.66 ;
      LAYER Metal6 ;
        RECT 181.66 12.00 182.32 12.66 ;
      LAYER Metal3 ;
        RECT 181.66 12.00 182.32 12.66 ;
      LAYER Metal4 ;
        RECT 181.66 12.00 182.32 12.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 224.98 12.00 225.64 12.66 ;
      LAYER Metal6 ;
        RECT 224.98 12.00 225.64 12.66 ;
      LAYER Metal3 ;
        RECT 224.98 12.00 225.64 12.66 ;
      LAYER Metal4 ;
        RECT 224.98 12.00 225.64 12.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 238.52 12.00 239.18 12.66 ;
      LAYER Metal6 ;
        RECT 238.52 12.00 239.18 12.66 ;
      LAYER Metal3 ;
        RECT 238.52 12.00 239.18 12.66 ;
      LAYER Metal4 ;
        RECT 238.52 12.00 239.18 12.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 246.26 12.00 246.92 12.66 ;
      LAYER Metal6 ;
        RECT 246.26 12.00 246.92 12.66 ;
      LAYER Metal3 ;
        RECT 246.26 12.00 246.92 12.66 ;
      LAYER Metal4 ;
        RECT 246.26 12.00 246.92 12.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 259.80 12.00 260.46 12.66 ;
      LAYER Metal6 ;
        RECT 259.80 12.00 260.46 12.66 ;
      LAYER Metal3 ;
        RECT 259.80 12.00 260.46 12.66 ;
      LAYER Metal4 ;
        RECT 259.80 12.00 260.46 12.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 32.70 12.00 33.36 12.66 ;
      LAYER Metal6 ;
        RECT 32.70 12.00 33.36 12.66 ;
      LAYER Metal3 ;
        RECT 32.70 12.00 33.36 12.66 ;
      LAYER Metal4 ;
        RECT 32.70 12.00 33.36 12.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 267.54 12.00 268.20 12.66 ;
      LAYER Metal6 ;
        RECT 267.54 12.00 268.20 12.66 ;
      LAYER Metal3 ;
        RECT 267.54 12.00 268.20 12.66 ;
      LAYER Metal4 ;
        RECT 267.54 12.00 268.20 12.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 281.08 12.00 281.74 12.66 ;
      LAYER Metal6 ;
        RECT 281.08 12.00 281.74 12.66 ;
      LAYER Metal3 ;
        RECT 281.08 12.00 281.74 12.66 ;
      LAYER Metal4 ;
        RECT 281.08 12.00 281.74 12.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 288.82 12.00 289.48 12.66 ;
      LAYER Metal6 ;
        RECT 288.82 12.00 289.48 12.66 ;
      LAYER Metal3 ;
        RECT 288.82 12.00 289.48 12.66 ;
      LAYER Metal4 ;
        RECT 288.82 12.00 289.48 12.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 302.36 12.00 303.02 12.66 ;
      LAYER Metal6 ;
        RECT 302.36 12.00 303.02 12.66 ;
      LAYER Metal3 ;
        RECT 302.36 12.00 303.02 12.66 ;
      LAYER Metal4 ;
        RECT 302.36 12.00 303.02 12.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 310.10 12.00 310.76 12.66 ;
      LAYER Metal6 ;
        RECT 310.10 12.00 310.76 12.66 ;
      LAYER Metal3 ;
        RECT 310.10 12.00 310.76 12.66 ;
      LAYER Metal4 ;
        RECT 310.10 12.00 310.76 12.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 323.64 12.00 324.30 12.66 ;
      LAYER Metal6 ;
        RECT 323.64 12.00 324.30 12.66 ;
      LAYER Metal3 ;
        RECT 323.64 12.00 324.30 12.66 ;
      LAYER Metal4 ;
        RECT 323.64 12.00 324.30 12.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 331.38 12.00 332.04 12.66 ;
      LAYER Metal6 ;
        RECT 331.38 12.00 332.04 12.66 ;
      LAYER Metal3 ;
        RECT 331.38 12.00 332.04 12.66 ;
      LAYER Metal4 ;
        RECT 331.38 12.00 332.04 12.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 344.92 12.00 345.58 12.66 ;
      LAYER Metal6 ;
        RECT 344.92 12.00 345.58 12.66 ;
      LAYER Metal3 ;
        RECT 344.92 12.00 345.58 12.66 ;
      LAYER Metal4 ;
        RECT 344.92 12.00 345.58 12.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 352.66 12.00 353.32 12.66 ;
      LAYER Metal6 ;
        RECT 352.66 12.00 353.32 12.66 ;
      LAYER Metal3 ;
        RECT 352.66 12.00 353.32 12.66 ;
      LAYER Metal4 ;
        RECT 352.66 12.00 353.32 12.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 366.20 12.00 366.86 12.66 ;
      LAYER Metal6 ;
        RECT 366.20 12.00 366.86 12.66 ;
      LAYER Metal3 ;
        RECT 366.20 12.00 366.86 12.66 ;
      LAYER Metal4 ;
        RECT 366.20 12.00 366.86 12.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 40.44 12.00 41.10 12.66 ;
      LAYER Metal6 ;
        RECT 40.44 12.00 41.10 12.66 ;
      LAYER Metal3 ;
        RECT 40.44 12.00 41.10 12.66 ;
      LAYER Metal4 ;
        RECT 40.44 12.00 41.10 12.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 373.94 12.00 374.60 12.66 ;
      LAYER Metal6 ;
        RECT 373.94 12.00 374.60 12.66 ;
      LAYER Metal3 ;
        RECT 373.94 12.00 374.60 12.66 ;
      LAYER Metal4 ;
        RECT 373.94 12.00 374.60 12.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 388.36 12.00 389.02 12.66 ;
      LAYER Metal6 ;
        RECT 388.36 12.00 389.02 12.66 ;
      LAYER Metal3 ;
        RECT 388.36 12.00 389.02 12.66 ;
      LAYER Metal4 ;
        RECT 388.36 12.00 389.02 12.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 53.98 12.00 54.64 12.66 ;
      LAYER Metal6 ;
        RECT 53.98 12.00 54.64 12.66 ;
      LAYER Metal3 ;
        RECT 53.98 12.00 54.64 12.66 ;
      LAYER Metal4 ;
        RECT 53.98 12.00 54.64 12.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 61.72 12.00 62.38 12.66 ;
      LAYER Metal6 ;
        RECT 61.72 12.00 62.38 12.66 ;
      LAYER Metal3 ;
        RECT 61.72 12.00 62.38 12.66 ;
      LAYER Metal4 ;
        RECT 61.72 12.00 62.38 12.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 75.26 12.00 75.92 12.66 ;
      LAYER Metal6 ;
        RECT 75.26 12.00 75.92 12.66 ;
      LAYER Metal3 ;
        RECT 75.26 12.00 75.92 12.66 ;
      LAYER Metal4 ;
        RECT 75.26 12.00 75.92 12.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 83.00 12.00 83.66 12.66 ;
      LAYER Metal6 ;
        RECT 83.00 12.00 83.66 12.66 ;
      LAYER Metal3 ;
        RECT 83.00 12.00 83.66 12.66 ;
      LAYER Metal4 ;
        RECT 83.00 12.00 83.66 12.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 96.54 12.00 97.20 12.66 ;
      LAYER Metal6 ;
        RECT 96.54 12.00 97.20 12.66 ;
      LAYER Metal3 ;
        RECT 96.54 12.00 97.20 12.66 ;
      LAYER Metal4 ;
        RECT 96.54 12.00 97.20 12.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 104.28 12.00 104.94 12.66 ;
      LAYER Metal6 ;
        RECT 104.28 12.00 104.94 12.66 ;
      LAYER Metal3 ;
        RECT 104.28 12.00 104.94 12.66 ;
      LAYER Metal4 ;
        RECT 104.28 12.00 104.94 12.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 117.82 12.00 118.48 12.66 ;
      LAYER Metal6 ;
        RECT 117.82 12.00 118.48 12.66 ;
      LAYER Metal3 ;
        RECT 117.82 12.00 118.48 12.66 ;
      LAYER Metal4 ;
        RECT 117.82 12.00 118.48 12.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 22.06 12.00 22.72 12.66 ;
      LAYER Metal6 ;
        RECT 22.06 12.00 22.72 12.66 ;
      LAYER Metal3 ;
        RECT 22.06 12.00 22.72 12.66 ;
      LAYER Metal4 ;
        RECT 22.06 12.00 22.72 12.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 128.46 12.00 129.12 12.66 ;
      LAYER Metal6 ;
        RECT 128.46 12.00 129.12 12.66 ;
      LAYER Metal3 ;
        RECT 128.46 12.00 129.12 12.66 ;
      LAYER Metal4 ;
        RECT 128.46 12.00 129.12 12.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 136.20 12.00 136.86 12.66 ;
      LAYER Metal6 ;
        RECT 136.20 12.00 136.86 12.66 ;
      LAYER Metal3 ;
        RECT 136.20 12.00 136.86 12.66 ;
      LAYER Metal4 ;
        RECT 136.20 12.00 136.86 12.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 149.74 12.00 150.40 12.66 ;
      LAYER Metal6 ;
        RECT 149.74 12.00 150.40 12.66 ;
      LAYER Metal3 ;
        RECT 149.74 12.00 150.40 12.66 ;
      LAYER Metal4 ;
        RECT 149.74 12.00 150.40 12.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 157.48 12.00 158.14 12.66 ;
      LAYER Metal6 ;
        RECT 157.48 12.00 158.14 12.66 ;
      LAYER Metal3 ;
        RECT 157.48 12.00 158.14 12.66 ;
      LAYER Metal4 ;
        RECT 157.48 12.00 158.14 12.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 171.02 12.00 171.68 12.66 ;
      LAYER Metal6 ;
        RECT 171.02 12.00 171.68 12.66 ;
      LAYER Metal3 ;
        RECT 171.02 12.00 171.68 12.66 ;
      LAYER Metal4 ;
        RECT 171.02 12.00 171.68 12.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.76 12.00 179.42 12.66 ;
      LAYER Metal6 ;
        RECT 178.76 12.00 179.42 12.66 ;
      LAYER Metal3 ;
        RECT 178.76 12.00 179.42 12.66 ;
      LAYER Metal4 ;
        RECT 178.76 12.00 179.42 12.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 227.88 12.00 228.54 12.66 ;
      LAYER Metal6 ;
        RECT 227.88 12.00 228.54 12.66 ;
      LAYER Metal3 ;
        RECT 227.88 12.00 228.54 12.66 ;
      LAYER Metal4 ;
        RECT 227.88 12.00 228.54 12.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 235.62 12.00 236.28 12.66 ;
      LAYER Metal6 ;
        RECT 235.62 12.00 236.28 12.66 ;
      LAYER Metal3 ;
        RECT 235.62 12.00 236.28 12.66 ;
      LAYER Metal4 ;
        RECT 235.62 12.00 236.28 12.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 249.16 12.00 249.82 12.66 ;
      LAYER Metal6 ;
        RECT 249.16 12.00 249.82 12.66 ;
      LAYER Metal3 ;
        RECT 249.16 12.00 249.82 12.66 ;
      LAYER Metal4 ;
        RECT 249.16 12.00 249.82 12.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 256.90 12.00 257.56 12.66 ;
      LAYER Metal6 ;
        RECT 256.90 12.00 257.56 12.66 ;
      LAYER Metal3 ;
        RECT 256.90 12.00 257.56 12.66 ;
      LAYER Metal4 ;
        RECT 256.90 12.00 257.56 12.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 29.80 12.00 30.46 12.66 ;
      LAYER Metal6 ;
        RECT 29.80 12.00 30.46 12.66 ;
      LAYER Metal3 ;
        RECT 29.80 12.00 30.46 12.66 ;
      LAYER Metal4 ;
        RECT 29.80 12.00 30.46 12.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 270.44 12.00 271.10 12.66 ;
      LAYER Metal6 ;
        RECT 270.44 12.00 271.10 12.66 ;
      LAYER Metal3 ;
        RECT 270.44 12.00 271.10 12.66 ;
      LAYER Metal4 ;
        RECT 270.44 12.00 271.10 12.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 278.18 12.00 278.84 12.66 ;
      LAYER Metal6 ;
        RECT 278.18 12.00 278.84 12.66 ;
      LAYER Metal3 ;
        RECT 278.18 12.00 278.84 12.66 ;
      LAYER Metal4 ;
        RECT 278.18 12.00 278.84 12.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.72 12.00 292.38 12.66 ;
      LAYER Metal6 ;
        RECT 291.72 12.00 292.38 12.66 ;
      LAYER Metal3 ;
        RECT 291.72 12.00 292.38 12.66 ;
      LAYER Metal4 ;
        RECT 291.72 12.00 292.38 12.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 299.46 12.00 300.12 12.66 ;
      LAYER Metal6 ;
        RECT 299.46 12.00 300.12 12.66 ;
      LAYER Metal3 ;
        RECT 299.46 12.00 300.12 12.66 ;
      LAYER Metal4 ;
        RECT 299.46 12.00 300.12 12.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 313.00 12.00 313.66 12.66 ;
      LAYER Metal6 ;
        RECT 313.00 12.00 313.66 12.66 ;
      LAYER Metal3 ;
        RECT 313.00 12.00 313.66 12.66 ;
      LAYER Metal4 ;
        RECT 313.00 12.00 313.66 12.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 320.74 12.00 321.40 12.66 ;
      LAYER Metal6 ;
        RECT 320.74 12.00 321.40 12.66 ;
      LAYER Metal3 ;
        RECT 320.74 12.00 321.40 12.66 ;
      LAYER Metal4 ;
        RECT 320.74 12.00 321.40 12.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 334.28 12.00 334.94 12.66 ;
      LAYER Metal6 ;
        RECT 334.28 12.00 334.94 12.66 ;
      LAYER Metal3 ;
        RECT 334.28 12.00 334.94 12.66 ;
      LAYER Metal4 ;
        RECT 334.28 12.00 334.94 12.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 342.02 12.00 342.68 12.66 ;
      LAYER Metal6 ;
        RECT 342.02 12.00 342.68 12.66 ;
      LAYER Metal3 ;
        RECT 342.02 12.00 342.68 12.66 ;
      LAYER Metal4 ;
        RECT 342.02 12.00 342.68 12.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 355.56 12.00 356.22 12.66 ;
      LAYER Metal6 ;
        RECT 355.56 12.00 356.22 12.66 ;
      LAYER Metal3 ;
        RECT 355.56 12.00 356.22 12.66 ;
      LAYER Metal4 ;
        RECT 355.56 12.00 356.22 12.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 363.30 12.00 363.96 12.66 ;
      LAYER Metal6 ;
        RECT 363.30 12.00 363.96 12.66 ;
      LAYER Metal3 ;
        RECT 363.30 12.00 363.96 12.66 ;
      LAYER Metal4 ;
        RECT 363.30 12.00 363.96 12.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 43.34 12.00 44.00 12.66 ;
      LAYER Metal6 ;
        RECT 43.34 12.00 44.00 12.66 ;
      LAYER Metal3 ;
        RECT 43.34 12.00 44.00 12.66 ;
      LAYER Metal4 ;
        RECT 43.34 12.00 44.00 12.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.84 12.00 377.50 12.66 ;
      LAYER Metal6 ;
        RECT 376.84 12.00 377.50 12.66 ;
      LAYER Metal3 ;
        RECT 376.84 12.00 377.50 12.66 ;
      LAYER Metal4 ;
        RECT 376.84 12.00 377.50 12.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.58 12.00 385.24 12.66 ;
      LAYER Metal6 ;
        RECT 384.58 12.00 385.24 12.66 ;
      LAYER Metal3 ;
        RECT 384.58 12.00 385.24 12.66 ;
      LAYER Metal4 ;
        RECT 384.58 12.00 385.24 12.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 51.08 12.00 51.74 12.66 ;
      LAYER Metal6 ;
        RECT 51.08 12.00 51.74 12.66 ;
      LAYER Metal3 ;
        RECT 51.08 12.00 51.74 12.66 ;
      LAYER Metal4 ;
        RECT 51.08 12.00 51.74 12.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.62 12.00 65.28 12.66 ;
      LAYER Metal6 ;
        RECT 64.62 12.00 65.28 12.66 ;
      LAYER Metal3 ;
        RECT 64.62 12.00 65.28 12.66 ;
      LAYER Metal4 ;
        RECT 64.62 12.00 65.28 12.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.36 12.00 73.02 12.66 ;
      LAYER Metal6 ;
        RECT 72.36 12.00 73.02 12.66 ;
      LAYER Metal3 ;
        RECT 72.36 12.00 73.02 12.66 ;
      LAYER Metal4 ;
        RECT 72.36 12.00 73.02 12.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.90 12.00 86.56 12.66 ;
      LAYER Metal6 ;
        RECT 85.90 12.00 86.56 12.66 ;
      LAYER Metal3 ;
        RECT 85.90 12.00 86.56 12.66 ;
      LAYER Metal4 ;
        RECT 85.90 12.00 86.56 12.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.64 12.00 94.30 12.66 ;
      LAYER Metal6 ;
        RECT 93.64 12.00 94.30 12.66 ;
      LAYER Metal3 ;
        RECT 93.64 12.00 94.30 12.66 ;
      LAYER Metal4 ;
        RECT 93.64 12.00 94.30 12.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.18 12.00 107.84 12.66 ;
      LAYER Metal6 ;
        RECT 107.18 12.00 107.84 12.66 ;
      LAYER Metal3 ;
        RECT 107.18 12.00 107.84 12.66 ;
      LAYER Metal4 ;
        RECT 107.18 12.00 107.84 12.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 114.92 12.00 115.58 12.66 ;
      LAYER Metal6 ;
        RECT 114.92 12.00 115.58 12.66 ;
      LAYER Metal3 ;
        RECT 114.92 12.00 115.58 12.66 ;
      LAYER Metal4 ;
        RECT 114.92 12.00 115.58 12.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 212.68 12.00 213.34 12.66 ;
      LAYER Metal6 ;
        RECT 212.68 12.00 213.34 12.66 ;
      LAYER Metal3 ;
        RECT 212.68 12.00 213.34 12.66 ;
      LAYER Metal4 ;
        RECT 212.68 12.00 213.34 12.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 193.96 12.00 194.62 12.66 ;
      LAYER Metal6 ;
        RECT 193.96 12.00 194.62 12.66 ;
      LAYER Metal3 ;
        RECT 193.96 12.00 194.62 12.66 ;
      LAYER Metal4 ;
        RECT 193.96 12.00 194.62 12.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 140.03 423.01 145.03 ;
        RECT 0.00 0.00 423.01 5.00 ;
      LAYER Metal2 ;
        RECT 418.01 0.00 423.01 145.03 ;
        RECT 0.00 0.00 5.00 145.03 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.60 134.44 417.42 139.44 ;
        RECT 5.60 5.60 417.42 10.60 ;
      LAYER Metal2 ;
        RECT 412.42 5.60 417.42 139.44 ;
        RECT 5.60 5.60 10.60 139.44 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12.00 12.00 411.02 132.97 ;
    LAYER Metal2 ;
      RECT 12.00 12.00 411.02 132.97 ;
    LAYER Metal3 ;
      RECT 12.00 12.00 411.02 132.97 ;
    LAYER Metal4 ;
      RECT 12.00 12.00 411.02 132.97 ;
    LAYER Metal5 ;
      RECT 12.00 12.00 411.02 132.97 ;
    LAYER Metal6 ;
      RECT 12.00 12.00 411.02 132.97 ;
  END
END MEM2


END LIBRARY

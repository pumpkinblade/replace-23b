VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


UNITS
  CAPACITANCE PICOFARADS 1 ;
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;


LAYER Metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.06 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0    0.06 
    WIDTH 0.1  0.1 
    WIDTH 0.75 0.25 
    WIDTH 1.5  0.45 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.15
    WIDTH 0.75  0.25
    WIDTH 1.5   0.45 ;
  SPACING 0.1 ENDOFLINE 0.1 WITHIN 0.035 ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.15
    WIDTH 0.75  0.25
    WIDTH 1.5   0.45 ;
  SPACING 0.1 ENDOFLINE 0.1 WITHIN 0.035 ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.15
    WIDTH 0.75  0.25
    WIDTH 1.5   0.45 ;
  SPACING 0.1 ENDOFLINE 0.1 WITHIN 0.035 ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.15
    WIDTH 0.75  0.25
    WIDTH 1.5   0.45 ;
  SPACING 0.1 ENDOFLINE 0.1 WITHIN 0.035 ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.15
    WIDTH 0.75  0.25
    WIDTH 1.5   0.45 ;
  SPACING 0.1 ENDOFLINE 0.1 WITHIN 0.035 ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.15
    WIDTH 0.75  0.25
    WIDTH 1.5   0.45 ;
  SPACING 0.1 ENDOFLINE 0.1 WITHIN 0.035 ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.15
    WIDTH 0.75  0.25
    WIDTH 1.5   0.45 ;
  SPACING 0.1 ENDOFLINE 0.1 WITHIN 0.035 ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.33 0.33 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.15
    WIDTH 0.75  0.25
    WIDTH 1.5   0.45 ;
  SPACING 0.1 ENDOFLINE 0.1 WITHIN 0.035 ;
END Metal9

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1C DEFAULT 
    LAYER Metal1 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER Metal1 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal2 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER Metal1 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA12_1C_V

VIA VIA23_1C DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER Metal2 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA23_1C_V

VIA VIA23_1ST_N DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.325000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1ST_N

VIA VIA23_1ST_S DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.325000 0.035000 0.065000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1ST_S

VIA VIA34_1C DEFAULT 
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER Metal3 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1C_V

VIA VIA34_1ST_E DEFAULT 
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.325000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1ST_E

VIA VIA34_1ST_W DEFAULT 
    LAYER Metal3 ;
        RECT -0.325000 -0.035000 0.065000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1ST_W

VIA VIA45_1C DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1C

VIA VIA45_1C_H DEFAULT 
    LAYER Metal4 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1C_H

VIA VIA45_1C_V DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA45_1C_V

VIA VIA45_1ST_N DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.325000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1ST_N

VIA VIA45_1ST_S DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.325000 0.035000 0.065000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1ST_S

VIA VIA5_0_VH DEFAULT 
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via5 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA5_0_VH

VIA VIA6_0_HV DEFAULT 
    LAYER Metal6 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
    LAYER Via6 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER Metal7 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
END VIA6_0_HV

VIA VIA7_0_VH DEFAULT 
    LAYER Metal7 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
    LAYER Via7 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER Metal8 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
END VIA7_0_VH

VIA VIA8_0_VH DEFAULT 
    LAYER Metal8 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
    LAYER Via8 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER Metal9 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
END VIA8_0_VH


SITE CoreSite
  CLASS CORE ;
  SIZE 0.2 BY 1.71 ;
END CoreSite

MACRO OAI2BB1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X4 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 0.59 0.175 1.22 ;
        RECT 0.06 0.98 0.175 1.22 ;
        RECT 0.335 1.16 0.395 1.44 ;
        RECT 0.51 0.57 0.63 0.65 ;
        RECT 0.745 1.16 0.805 1.44 ;
        RECT 0.115 0.59 1.145 0.65 ;
        RECT 1.165 1.16 1.225 1.44 ;
        RECT 1.095 0.57 1.36 0.63 ;
        RECT 0.06 1.16 1.635 1.22 ;
        RECT 1.575 1.16 1.635 1.44 ;
    END
  END Y
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 0.625 1.965 0.705 ;
        RECT 1.885 0.625 1.965 0.9 ;
        RECT 1.885 0.82 2.1 0.9 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.36 0.76 2.44 1.06 ;
        RECT 2.36 0.98 2.54 1.06 ;
        RECT 2.46 0.98 2.54 1.16 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.75 0.54 0.92 ;
        RECT 0.275 0.75 1.695 0.81 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END OAI2BB1X4

MACRO OA22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.67 1.5 1.395 ;
        RECT 1.46 0.57 1.54 0.73 ;
        RECT 1.46 0.57 1.615 0.63 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.98 1.08 1.17 ;
        RECT 1 0.98 1.34 1.06 ;
        RECT 1.26 0.98 1.34 1.11 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.675 0.54 1.175 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.675 0.34 1.175 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.675 0.74 1.175 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END OA22X2

MACRO NAND3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X8 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.315 1.195 0.375 1.46 ;
        RECT 0.76 1.21 0.82 1.33 ;
        RECT 1.17 1.21 1.23 1.33 ;
        RECT 1.58 1.06 1.64 1.46 ;
        RECT 2.025 1.21 2.085 1.33 ;
        RECT 2.44 1.21 2.5 1.33 ;
        RECT 2.85 1.21 2.91 1.33 ;
        RECT 3.26 1.21 3.32 1.33 ;
        RECT 3.705 1.06 3.765 1.46 ;
        RECT 0.315 1.21 4.175 1.27 ;
        RECT 4.115 1.015 4.175 1.46 ;
        RECT 4.46 0.98 4.625 1.11 ;
        RECT 4.115 1.05 4.625 1.11 ;
        RECT 0.775 0.405 4.625 0.465 ;
        RECT 4.565 0.405 4.625 1.46 ;
        RECT 4.525 0.98 4.625 1.46 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.28 0.79 0.34 1.095 ;
        RECT 0.28 1.035 0.535 1.095 ;
        RECT 1.28 0.885 1.34 1.11 ;
        RECT 0.475 1.05 1.34 1.11 ;
        RECT 1.28 0.885 1.4 0.96 ;
        RECT 1.28 0.9 1.8 0.96 ;
        RECT 1.74 0.9 1.8 1.11 ;
        RECT 2.55 0.885 2.67 0.945 ;
        RECT 2.61 0.885 2.67 1.11 ;
        RECT 3.545 0.9 3.605 1.11 ;
        RECT 1.74 1.05 3.605 1.11 ;
        RECT 3.545 0.9 3.79 0.96 ;
        RECT 3.73 0.885 3.86 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 0.875 0.695 0.935 ;
        RECT 1.04 0.725 1.1 0.95 ;
        RECT 0.635 0.89 1.1 0.95 ;
        RECT 1.04 0.725 1.56 0.785 ;
        RECT 1.5 0.74 1.96 0.8 ;
        RECT 1.9 0.74 1.96 0.95 ;
        RECT 2.28 0.74 2.34 0.95 ;
        RECT 1.9 0.89 2.34 0.95 ;
        RECT 2.28 0.74 2.4 0.8 ;
        RECT 2.34 0.725 2.83 0.785 ;
        RECT 2.77 0.74 3.03 0.8 ;
        RECT 2.97 0.74 3.03 0.95 ;
        RECT 3.385 0.74 3.445 0.95 ;
        RECT 2.97 0.89 3.445 0.95 ;
        RECT 3.385 0.74 3.63 0.8 ;
        RECT 3.51 0.725 4.245 0.785 ;
        RECT 4.035 0.725 4.245 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 0.79 ;
        RECT 0.795 0.73 0.94 0.79 ;
        RECT 2.06 0.565 2.12 0.79 ;
        RECT 2.06 0.73 2.18 0.79 ;
        RECT 3.225 0.565 3.285 0.79 ;
        RECT 3.165 0.73 3.285 0.79 ;
        RECT 0.88 0.565 4.405 0.625 ;
        RECT 4.345 0.565 4.405 0.8 ;
        RECT 4.345 0.74 4.465 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END NAND3X8

MACRO SDFFRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX4 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.66 0.485 6.72 1.34 ;
        RECT 6.66 0.79 6.74 1.34 ;
        RECT 6.66 0.95 6.76 1.34 ;
        RECT 6.66 0.95 7.17 1.01 ;
        RECT 7.11 0.95 7.17 1.34 ;
        RECT 6.6 0.485 7.19 0.545 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.86 0.485 5.92 1.34 ;
        RECT 5.86 0.79 5.94 1.34 ;
        RECT 5.66 0.485 6.25 0.545 ;
        RECT 5.86 0.95 6.35 1.01 ;
        RECT 6.29 0.95 6.35 1.34 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.635 0.625 3.765 0.705 ;
        RECT 3.705 0.295 3.765 0.865 ;
        RECT 3.225 0.805 3.765 0.865 ;
        RECT 3.705 0.295 4.47 0.355 ;
        RECT 4.41 0.295 4.47 0.45 ;
        RECT 4.41 0.39 4.785 0.45 ;
        RECT 4.725 0.39 4.785 0.705 ;
        RECT 4.725 0.64 5.41 0.705 ;
        RECT 4.665 0.645 5.41 0.705 ;
        RECT 5.35 0.64 5.41 0.76 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.6 1.54 1.1 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.6 1.34 1.1 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.74 0.54 1.1 ;
        RECT 0.46 0.79 0.68 1.1 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.54 0.255 0.6 0.64 ;
        RECT 0.28 0.58 0.695 0.64 ;
        RECT 0.635 0.625 0.755 0.685 ;
        RECT 0.54 0.255 1.16 0.315 ;
        RECT 1.1 0.255 1.16 1.1 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.8 0.06 ;
    END
  END VSS
END SDFFRX4

MACRO TLATSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRX1 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 0.73 ;
        RECT 0.88 0.41 0.94 1.07 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.305 0.54 ;
        RECT 0.225 0.41 0.305 1.29 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.39 0.785 3.47 1.155 ;
        RECT 3.26 0.845 3.47 1.155 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.025 0.785 2.105 0.96 ;
        RECT 2.025 0.815 2.43 0.96 ;
    END
  END RN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 0.815 1.68 1.23 ;
        RECT 1.6 0.815 1.765 0.895 ;
    END
  END G
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.2 0.84 1.34 0.92 ;
        RECT 1.26 0.65 1.34 1.09 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END TLATSRX1

MACRO OAI2BB1X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.18 0.54 ;
        RECT 0.12 0.4 0.18 0.85 ;
        RECT 0.12 0.79 0.34 0.85 ;
        RECT 0.28 0.79 0.34 1.34 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.64 0.52 1.06 ;
        RECT 0.46 0.98 0.54 1.12 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.64 0.72 1.12 ;
        RECT 0.64 0.78 0.74 1.12 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.67 1.08 1.06 ;
        RECT 1.06 0.98 1.14 1.11 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OAI2BB1X1

MACRO DLY4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY4X1 0 0 ;
  SIZE 5.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.54 0.515 1.29 ;
        RECT 0.435 0.625 0.565 0.705 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.46 0.69 5.54 1.19 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.8 0.06 ;
    END
  END VSS
END DLY4X1

MACRO ADDFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.745 0.415 4.805 0.555 ;
        RECT 4.745 1 4.805 1.39 ;
        RECT 4.745 0.495 5.285 0.555 ;
        RECT 5.155 1 5.215 1.39 ;
        RECT 5.165 0.415 5.225 0.555 ;
        RECT 5.225 0.495 5.285 1.06 ;
        RECT 4.745 1 5.285 1.06 ;
        RECT 5.225 0.6 5.34 0.73 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.28 0.6 0.34 0.98 ;
        RECT 0.34 0.52 0.4 0.66 ;
        RECT 0.34 0.92 0.4 1.295 ;
        RECT 0.28 0.92 0.82 0.98 ;
        RECT 0.76 0.52 0.82 0.66 ;
        RECT 0.26 0.6 0.82 0.66 ;
        RECT 0.76 0.92 0.82 1.295 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 0.79 2.525 0.85 ;
        RECT 2.26 0.79 2.525 0.94 ;
        RECT 2.26 0.88 3.235 0.94 ;
        RECT 3.175 0.82 4.325 0.88 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.54 0.63 1.6 0.75 ;
        RECT 1.54 0.63 2.685 0.69 ;
        RECT 2.625 0.63 2.685 0.78 ;
        RECT 2.625 0.72 3.075 0.78 ;
        RECT 3.015 0.66 4.485 0.72 ;
        RECT 4.235 0.625 4.485 0.72 ;
        RECT 4.425 0.625 4.485 0.745 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.435 2.365 0.53 ;
        RECT 2.235 0.47 2.825 0.53 ;
        RECT 2.795 0.5 2.915 0.62 ;
        RECT 2.765 0.5 4.015 0.56 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END ADDFX4

MACRO CLKAND2X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X12 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.305 0.35 2.365 0.655 ;
        RECT 2.395 0.915 2.455 1.37 ;
        RECT 2.715 0.35 2.775 0.655 ;
        RECT 2.805 0.915 2.865 1.37 ;
        RECT 3.125 0.35 3.185 0.655 ;
        RECT 3.215 0.915 3.275 1.37 ;
        RECT 3.535 0.35 3.595 0.655 ;
        RECT 3.625 0.915 3.685 1.37 ;
        RECT 3.945 0.35 4.005 0.655 ;
        RECT 2.395 0.915 4.14 0.975 ;
        RECT 2.305 0.595 4.12 0.655 ;
        RECT 4.06 0.595 4.12 1.37 ;
        RECT 4.06 0.79 4.14 1.37 ;
        RECT 4.035 0.915 4.14 1.37 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.89 0.72 1.01 ;
        RECT 1.19 0.89 1.25 1.01 ;
        RECT 1.835 0.815 1.965 1.01 ;
        RECT 0.66 0.95 1.965 1.01 ;
        RECT 1.835 0.815 2.045 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 0.79 0.54 0.85 ;
        RECT 0.46 0.79 0.54 0.92 ;
        RECT 0.965 0.73 1.085 0.8 ;
        RECT 0.48 0.73 1.64 0.79 ;
        RECT 1.58 0.73 1.64 0.85 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END CLKAND2X12

MACRO MXI3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3XL 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.52 3.34 1.02 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 0.74 2.995 1.085 ;
        RECT 2.915 0.79 3.15 1.085 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 0.815 2.165 1.02 ;
        RECT 2.035 0.94 2.565 1.02 ;
    END
  END S1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.345 0.845 1.54 1.135 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.425 0.815 0.925 0.895 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.965 0.325 1.085 ;
        RECT 0.235 1.005 0.365 1.085 ;
        RECT 0.245 0.995 0.9 1.075 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END MXI3XL

MACRO NAND3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X6 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1.18 0.45 1.3 ;
        RECT 0.775 0.32 0.835 0.6 ;
        RECT 0.8 1.18 0.86 1.3 ;
        RECT 1.21 1.18 1.27 1.3 ;
        RECT 1.62 1.18 1.68 1.3 ;
        RECT 0.775 0.32 2.025 0.38 ;
        RECT 1.965 0.32 2.025 0.6 ;
        RECT 2.17 1.18 2.23 1.3 ;
        RECT 2.605 1.07 2.665 1.43 ;
        RECT 3.015 1.18 3.075 1.3 ;
        RECT 1.965 0.43 3.465 0.49 ;
        RECT 3.405 0.32 3.465 0.6 ;
        RECT 3.425 1.18 3.485 1.3 ;
        RECT 3.835 1.18 3.895 1.43 ;
        RECT 3.405 0.54 4.14 0.6 ;
        RECT 4.06 0.98 4.14 1.24 ;
        RECT 4.08 0.54 4.14 1.24 ;
        RECT 0.39 1.18 4.14 1.24 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.815 0.405 0.895 ;
        RECT 0.345 0.815 0.405 1.08 ;
        RECT 1.425 0.91 1.545 1.08 ;
        RECT 2.445 0.91 2.505 1.08 ;
        RECT 0.345 1.02 2.505 1.08 ;
        RECT 2.445 0.91 2.985 0.97 ;
        RECT 2.925 0.91 2.985 1.08 ;
        RECT 3.9 0.76 3.96 1.08 ;
        RECT 2.925 1.02 3.96 1.08 ;
        RECT 3.9 0.76 3.97 0.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.505 0.86 1.165 0.92 ;
        RECT 1.105 0.805 1.325 0.865 ;
        RECT 1.265 0.75 1.705 0.81 ;
        RECT 1.645 0.75 1.705 0.92 ;
        RECT 2.285 0.75 2.345 0.92 ;
        RECT 1.645 0.86 2.345 0.92 ;
        RECT 2.285 0.75 3.145 0.81 ;
        RECT 3.085 0.75 3.145 0.92 ;
        RECT 3.66 0.79 3.74 0.92 ;
        RECT 3.085 0.86 3.795 0.92 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 0.7 1.005 0.76 ;
        RECT 0.945 0.625 1.165 0.705 ;
        RECT 1.105 0.59 1.865 0.65 ;
        RECT 1.805 0.59 1.865 0.76 ;
        RECT 2.125 0.59 2.185 0.76 ;
        RECT 1.805 0.7 2.185 0.76 ;
        RECT 2.125 0.59 3.305 0.65 ;
        RECT 3.245 0.59 3.305 0.76 ;
        RECT 3.245 0.7 3.415 0.76 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.2 0.06 ;
    END
  END VSS
END NAND3X6

MACRO SDFFRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX2 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.055 0.49 1.135 0.99 ;
        RECT 1.055 0.6 1.14 0.73 ;
        RECT 1.055 0.91 1.175 0.99 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.49 0.73 0.99 ;
        RECT 0.56 0.91 0.73 0.99 ;
        RECT 0.65 0.6 0.74 0.73 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.635 0.6 5.715 0.88 ;
        RECT 5.635 0.6 6.14 0.68 ;
        RECT 6.06 0.6 6.14 0.73 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.815 0.78 5.895 1.085 ;
        RECT 5.635 1.005 5.895 1.085 ;
        RECT 5.815 0.78 5.935 0.86 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.79 5.14 1.025 ;
        RECT 5.135 0.6 5.215 0.87 ;
    END
  END SI
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.385 0.84 2.52 0.9 ;
        RECT 2.46 0.84 2.52 1.11 ;
        RECT 2.46 0.98 2.54 1.11 ;
        RECT 2.46 1.05 2.84 1.11 ;
        RECT 2.78 1.05 2.84 1.44 ;
        RECT 2.78 1.38 3.77 1.44 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.57 1.515 0.945 ;
        RECT 1.435 0.57 1.64 0.705 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END SDFFRX2

MACRO MX3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X1 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.08 0.41 0.14 0.825 ;
        RECT 0.13 0.385 0.19 0.505 ;
        RECT 0.13 0.765 0.19 1.345 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.08 0.965 2.16 1.085 ;
        RECT 2.08 1.005 2.765 1.085 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.775 2.34 0.905 ;
        RECT 2.26 0.775 2.71 0.855 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.6 1.54 0.73 ;
        RECT 1.46 0.65 1.66 0.73 ;
        RECT 1.58 0.65 1.66 0.98 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.48 1.34 0.98 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.625 0.54 1.125 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END MX3X1

MACRO SDFFSRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX1 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.51 0.14 0.73 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.11 0.67 0.17 1.29 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.825 0.645 6.885 0.905 ;
        RECT 7.39 0.625 7.565 0.705 ;
        RECT 6.825 0.645 7.565 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.235 0.805 7.34 0.98 ;
        RECT 7.205 0.81 7.34 0.98 ;
        RECT 7.205 0.815 7.61 0.895 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.435 0.54 6.565 0.91 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.85 0.815 6.165 0.91 ;
        RECT 5.85 0.815 6.335 0.895 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.79 1.54 0.92 ;
        RECT 1.48 0.79 1.54 1.005 ;
        RECT 1.48 0.945 2.46 1.005 ;
        RECT 2.4 0.945 2.46 1.355 ;
        RECT 3.2 1.16 3.26 1.355 ;
        RECT 2.4 1.295 3.26 1.355 ;
        RECT 3.2 1.16 3.64 1.22 ;
        RECT 3.58 1.16 3.64 1.385 ;
        RECT 3.58 1.325 4.28 1.385 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 0.655 1.105 0.91 ;
        RECT 1.025 0.79 1.34 0.91 ;
        RECT 1.26 0.79 1.34 0.92 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.8 0.06 ;
    END
  END VSS
END SDFFSRHQX1

MACRO TLATNTSCAX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX16 0 0 ;
  SIZE 7.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.615 0.5 4.675 0.62 ;
        RECT 4.66 0.56 4.72 1.405 ;
        RECT 4.66 0.79 4.74 0.92 ;
        RECT 4.995 0.57 5.115 0.63 ;
        RECT 5.07 0.815 5.13 1.405 ;
        RECT 5.07 0.585 5.495 0.645 ;
        RECT 5.435 0.525 5.495 0.875 ;
        RECT 5.48 0.815 5.54 1.405 ;
        RECT 5.815 0.57 5.935 0.63 ;
        RECT 5.89 0.815 5.95 1.405 ;
        RECT 5.89 0.585 6.315 0.645 ;
        RECT 6.255 0.525 6.315 0.875 ;
        RECT 6.3 0.815 6.36 1.405 ;
        RECT 6.635 0.57 6.755 0.63 ;
        RECT 6.71 0.815 6.77 1.405 ;
        RECT 6.71 0.585 7.135 0.645 ;
        RECT 4.66 0.815 7.18 0.875 ;
        RECT 7.075 0.525 7.135 0.875 ;
        RECT 7.12 0.815 7.18 1.405 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.74 0.95 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.45 0.54 0.95 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.060 0.54 0.14 0.95 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.6 0.06 ;
    END
  END VSS
END TLATNTSCAX16

MACRO OAI33XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.965 1.185 1.025 1.37 ;
        RECT 1.14 0.29 1.26 0.35 ;
        RECT 1.2 0.29 1.26 0.485 ;
        RECT 1.595 0.26 1.74 0.485 ;
        RECT 1.2 0.425 1.74 0.485 ;
        RECT 1.66 0.98 1.74 1.245 ;
        RECT 1.68 0.26 1.74 1.245 ;
        RECT 0.965 1.185 1.74 1.245 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.745 0.54 1.245 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.775 0.94 1.085 ;
        RECT 0.86 1.005 1.13 1.085 ;
    END
  END B2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.06 0.65 0.32 0.73 ;
        RECT 0.22 0.65 0.32 0.92 ;
    END
  END A0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.79 0.74 1.29 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.585 1.34 1.085 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.585 1.52 0.705 ;
        RECT 1.46 0.6 1.54 1.065 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OAI33XL

MACRO TLATSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRX4 0 0 ;
  SIZE 7.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.465 3.72 1.055 ;
        RECT 3.66 0.79 3.74 1.055 ;
        RECT 4.1 0.675 4.16 1.055 ;
        RECT 3.6 0.995 4.22 1.055 ;
        RECT 4.36 0.465 4.42 0.735 ;
        RECT 4.1 0.675 4.42 0.735 ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.775 0.815 5.52 0.895 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.735 0.78 ;
        RECT 0.66 0.6 0.74 0.73 ;
        RECT 0.94 0.305 1 0.66 ;
        RECT 0.66 0.6 1 0.66 ;
        RECT 0.94 0.305 1.32 0.365 ;
        RECT 1.26 0.305 1.32 0.605 ;
        RECT 1.58 0.305 1.64 0.605 ;
        RECT 1.26 0.545 1.64 0.605 ;
        RECT 1.58 0.305 1.96 0.365 ;
        RECT 1.9 0.305 1.96 0.605 ;
        RECT 2.22 0.305 2.28 0.605 ;
        RECT 1.9 0.545 2.28 0.605 ;
        RECT 2.22 0.305 2.6 0.365 ;
        RECT 2.54 0.305 2.6 0.605 ;
        RECT 2.86 0.305 2.92 0.605 ;
        RECT 2.54 0.545 2.92 0.605 ;
        RECT 2.86 0.305 3.24 0.365 ;
        RECT 3.18 0.305 3.24 0.605 ;
        RECT 3.5 0.305 3.56 0.605 ;
        RECT 3.18 0.545 3.56 0.605 ;
        RECT 3.5 0.305 3.88 0.365 ;
        RECT 3.82 0.305 3.88 0.575 ;
        RECT 4.2 0.305 4.26 0.575 ;
        RECT 3.82 0.515 4.26 0.575 ;
        RECT 4.2 0.305 4.58 0.365 ;
        RECT 4.52 0.305 4.58 0.555 ;
        RECT 4.9 0.305 4.96 0.555 ;
        RECT 4.52 0.495 4.96 0.555 ;
        RECT 4.9 0.305 5.395 0.365 ;
        RECT 5.335 0.35 5.775 0.41 ;
        RECT 5.715 0.31 5.835 0.37 ;
    END
  END RN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.685 0.4 0.895 ;
        RECT 0.03 0.795 0.4 0.895 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.82 0.66 6.9 0.91 ;
        RECT 6.82 0.79 7.14 0.91 ;
        RECT 7.06 0.79 7.14 0.92 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.1 0.465 1.16 1.055 ;
        RECT 1.1 0.79 1.34 1.055 ;
        RECT 1.74 0.465 1.8 1.055 ;
        RECT 1.07 0.995 1.8 1.055 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.6 0.06 ;
    END
  END VSS
END TLATSRX4

MACRO DFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX4 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.1 0.815 4.6 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.43 0.34 0.93 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.545 0.57 0.74 0.63 ;
        RECT 0.66 0.57 0.74 0.73 ;
        RECT 0.68 0.57 0.74 1.29 ;
        RECT 0.66 0.67 1.105 0.73 ;
        RECT 1.045 0.54 1.105 0.99 ;
        RECT 1.09 0.93 1.15 1.29 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END DFFHQX4

MACRO AOI221X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X2 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.79 1.14 0.92 ;
        RECT 1.08 0.45 1.14 1.055 ;
        RECT 0.605 0.45 2.17 0.51 ;
        RECT 1.08 0.995 2.28 1.055 ;
        RECT 2.22 0.995 2.28 1.135 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.815 1.935 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.765 0.74 1.065 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.365 0.715 ;
        RECT 0.285 0.61 0.96 0.69 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.625 1.765 0.715 ;
        RECT 1.24 0.635 1.935 0.715 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.065 0.815 2.565 0.895 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END AOI221X2

MACRO ADDFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX2 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.255 0.42 4.315 1.09 ;
        RECT 4.255 0.6 4.34 0.73 ;
        RECT 4.225 1.03 4.345 1.09 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.06 0.79 0.335 0.85 ;
        RECT 0.275 0.54 0.335 1.31 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.19 0.81 1.47 0.87 ;
        RECT 2.06 0.82 2.14 1.11 ;
        RECT 1.425 0.82 3.735 0.88 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.97 0.685 1.09 0.745 ;
        RECT 1.03 0.65 1.57 0.71 ;
        RECT 1.53 0.66 3.965 0.72 ;
        RECT 3.835 0.66 3.965 0.895 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.435 1.765 0.56 ;
        RECT 1.635 0.5 3.515 0.56 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END ADDFX2

MACRO AOI22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 0.255 0.74 0.92 ;
        RECT 0.66 0.79 0.74 0.92 ;
        RECT 0.66 0.86 0.96 0.92 ;
        RECT 0.9 0.86 0.96 1.175 ;
        RECT 0.905 1.115 0.965 1.235 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.45 0.34 0.95 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.45 1.14 0.95 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 0.25 0.92 0.73 ;
        RECT 0.84 0.6 0.94 0.73 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.54 0.35 ;
        RECT 0.48 0.29 0.56 0.7 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END AOI22XL

MACRO NAND3BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.15 0.335 0.21 1.085 ;
        RECT 0.15 1.005 0.43 1.085 ;
        RECT 0.37 1.005 0.43 1.345 ;
        RECT 0.15 0.335 0.825 0.395 ;
        RECT 0.79 1.065 0.85 1.345 ;
        RECT 0.37 1.065 1.26 1.125 ;
        RECT 1.2 1.02 1.26 1.345 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.53 0.815 0.96 0.895 ;
        RECT 0.88 0.815 0.96 0.965 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.655 1.13 0.715 ;
        RECT 1.06 0.715 1.14 0.92 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.785 1.54 1.125 ;
        RECT 1.49 0.655 1.57 0.92 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END NAND3BX2

MACRO SDFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRXL 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.45 0.94 1.21 ;
        RECT 0.86 0.45 1.02 0.57 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.305 0.73 ;
        RECT 0.225 0.54 0.305 1.02 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.035 0.57 6.21 0.805 ;
        RECT 5.865 0.725 6.21 0.805 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.465 0.625 5.545 0.905 ;
        RECT 5.465 0.625 5.765 0.705 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.235 0.625 5.365 1.075 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.79 4.14 0.965 ;
        RECT 4.11 0.515 4.19 0.91 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.25 0.835 1.365 1.085 ;
        RECT 1.04 1.005 1.365 1.085 ;
        RECT 1.25 0.835 1.37 0.915 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END SDFFTRXL

MACRO OR3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X2 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.93 0.91 0.99 1.3 ;
        RECT 1.025 0.37 1.085 0.97 ;
        RECT 0.93 0.91 1.085 0.97 ;
        RECT 1.26 0.6 1.34 0.73 ;
        RECT 1.025 0.67 1.34 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 0.625 0.745 1.065 ;
        RECT 0.625 0.625 0.765 0.705 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.635 0.34 0.92 ;
        RECT 0.285 0.79 0.365 1.11 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.61 0.14 1.11 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END OR3X2

MACRO CLKBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX2 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.365 0.73 ;
        RECT 0.305 0.555 0.365 0.925 ;
        RECT 0.35 0.495 0.41 0.615 ;
        RECT 0.35 0.865 0.41 1.32 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.76 0.765 1.085 ;
        RECT 0.51 1.005 0.765 1.085 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END CLKBUFX2

MACRO TLATX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATX1 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.045 0.54 3.165 0.705 ;
        RECT 3.035 0.625 3.165 0.705 ;
        RECT 3.07 0.54 3.165 1.325 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.6 2.34 0.73 ;
        RECT 2.28 0.54 2.34 1.415 ;
    END
  END QN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.78 1.94 1.28 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.62 0.54 1.025 ;
        RECT 0.46 0.725 0.635 1.025 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END TLATX1

MACRO DFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX2 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.98 3.34 1.11 ;
        RECT 3.28 0.92 3.34 1.465 ;
        RECT 3.315 0.54 3.375 0.98 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.745 0.805 0.965 1.085 ;
        RECT 0.745 0.805 1.045 0.885 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.54 0.14 0.73 ;
        RECT 0.06 0.65 0.285 0.73 ;
        RECT 0.205 0.65 0.285 0.895 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END DFFHQX2

MACRO MXI4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4XL 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.215 0.73 ;
        RECT 0.135 0.54 0.215 1.02 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.435 0.815 3.935 0.895 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.435 0.995 3.89 1.085 ;
        RECT 3.485 0.995 3.89 1.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.775 0.745 2.855 1.085 ;
        RECT 2.775 1.005 3.015 1.085 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.3 0.88 2.565 1.085 ;
        RECT 2.3 0.88 2.675 0.96 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 0.625 1.765 0.705 ;
        RECT 1.685 0.625 1.765 0.985 ;
        RECT 1.685 0.905 1.82 0.985 ;
    END
  END D
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.48 0.27 0.54 0.83 ;
        RECT 0.48 0.71 0.545 0.83 ;
        RECT 1.06 0.245 1.18 0.33 ;
        RECT 0.48 0.27 1.39 0.33 ;
        RECT 1.33 0.27 1.39 0.96 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.2 0.06 ;
    END
  END VSS
END MXI4XL

MACRO AOI2BB2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X2 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.405 0.445 1.67 0.505 ;
        RECT 1.86 0.79 1.94 0.92 ;
        RECT 1.88 0.465 1.94 1.055 ;
        RECT 2.1 0.995 2.16 1.135 ;
        RECT 1.61 0.465 2.335 0.525 ;
        RECT 2.275 0.445 2.395 0.505 ;
        RECT 1.88 0.995 2.57 1.055 ;
        RECT 2.51 0.995 2.57 1.135 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.075 0.805 2.565 0.895 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.04 0.625 2.63 0.705 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.54 1.1 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.46 0.34 0.96 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END AOI2BB2X2

MACRO SEDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX2 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.86 0.6 5.065 0.73 ;
        RECT 4.985 0.52 5.065 1.02 ;
        RECT 4.985 0.52 5.19 0.6 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.535 0.885 4.615 1.02 ;
        RECT 4.6 0.52 4.68 0.99 ;
        RECT 4.535 0.885 4.685 0.99 ;
        RECT 4.6 0.52 4.72 0.6 ;
        RECT 4.6 0.79 4.74 0.92 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.835 0.615 7.955 1.065 ;
        RECT 7.835 0.815 7.965 1.065 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.495 0.775 7.575 0.895 ;
        RECT 7.035 0.815 7.575 0.895 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.76 0.815 6.025 1.13 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.68 4.34 1.18 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.19 0.805 0.67 0.895 ;
        RECT 0.19 0.815 0.68 0.895 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.435 0.705 ;
        RECT 0.635 0.3 0.695 0.705 ;
        RECT 0.235 0.645 0.84 0.705 ;
        RECT 0.635 0.3 1.16 0.36 ;
        RECT 1.1 0.3 1.16 0.85 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.2 0.06 ;
    END
  END VSS
END SEDFFTRX2

MACRO SDFFNSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX2 0 0 ;
  SIZE 8.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.835 0.625 7.965 0.705 ;
        RECT 7.885 0.535 7.965 0.99 ;
        RECT 7.91 0.495 7.99 0.615 ;
        RECT 7.885 0.91 8.02 0.99 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.98 7.465 1.11 ;
        RECT 7.405 0.495 7.465 1.41 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.46 0.42 0.64 0.54 ;
        RECT 0.195 0.46 0.64 0.54 ;
        RECT 0.56 0.42 0.64 0.545 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.33 3.34 0.705 ;
        RECT 3.26 0.625 3.465 0.705 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.65 1.14 1.15 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.38 0.64 0.46 1.02 ;
        RECT 0.26 0.79 0.46 1.02 ;
    END
  END SI
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.06 0.69 7.14 1.19 ;
    END
  END RN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.335 0.585 1.415 0.895 ;
        RECT 1.335 0.815 1.605 0.895 ;
    END
  END CKN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.6 0.06 ;
    END
  END VSS
END SDFFNSRX2

MACRO INVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX8 0 0 ;
  SIZE 1.80 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.485 0.72 1.565 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.72 0.15 0.87 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.80 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.80 0.06 ;
    END
  END VSS
END INVX8

MACRO AOI33X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.795 0.38 0.855 0.5 ;
        RECT 1 1.2 1.06 1.32 ;
        RECT 0.795 0.44 1.52 0.5 ;
        RECT 1 1.2 1.52 1.26 ;
        RECT 1.46 0.44 1.52 1.48 ;
        RECT 1.46 0.98 1.54 1.11 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.49 0.34 0.99 ;
    END
  END A0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 1.1 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.79 1.14 1.085 ;
        RECT 1.075 0.6 1.155 0.87 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.6 1.34 1.1 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.23 0.54 0.73 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 1.1 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END AOI33X1

MACRO OR4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.385 0.99 1.445 1.36 ;
        RECT 1.44 0.405 1.5 0.545 ;
        RECT 1.385 0.99 1.94 1.05 ;
        RECT 1.795 0.99 1.855 1.36 ;
        RECT 1.85 0.405 1.94 0.545 ;
        RECT 1.44 0.485 1.94 0.545 ;
        RECT 1.88 0.405 1.94 1.3 ;
        RECT 1.795 0.99 1.94 1.3 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.79 0.74 1.14 ;
        RECT 0.665 0.645 0.745 0.92 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.645 0.56 1.125 ;
        RECT 0.46 0.8 0.56 1.125 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.485 1.34 0.73 ;
        RECT 1.005 0.65 1.34 0.73 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END OR4X4

MACRO DFFNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX1 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.955 0.995 1.11 ;
        RECT 0.89 0.475 0.95 1.11 ;
        RECT 0.935 0.955 0.995 1.345 ;
        RECT 0.94 0.435 1 0.555 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.325 0.54 ;
        RECT 0.245 0.41 0.325 1.29 ;
    END
  END QN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.06 0.52 6.14 1.02 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.445 0.46 5.525 0.945 ;
        RECT 5.445 0.46 5.54 0.815 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.005 0.77 2.125 0.83 ;
        RECT 2.035 1.005 2.165 1.085 ;
        RECT 2.06 0.77 2.125 1.085 ;
        RECT 2.105 1.005 2.165 1.23 ;
        RECT 2.105 1.17 3.165 1.23 ;
        RECT 3.105 1.185 4.015 1.245 ;
        RECT 3.955 1.185 4.015 1.465 ;
        RECT 3.955 1.405 4.47 1.465 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.095 0.815 1.34 1.125 ;
        RECT 1.095 0.815 1.365 0.895 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END DFFNSRX1

MACRO NAND3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.055 0.43 1.335 ;
        RECT 0.78 1.055 0.84 1.335 ;
        RECT 1.19 1.055 1.25 1.335 ;
        RECT 0.795 0.335 1.565 0.395 ;
        RECT 1.435 1.005 1.565 1.115 ;
        RECT 1.505 0.335 1.565 1.115 ;
        RECT 0.36 1.055 1.565 1.115 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.52 0.815 0.765 0.955 ;
        RECT 0.52 0.815 0.96 0.895 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.655 1.14 0.715 ;
        RECT 1.06 0.655 1.14 0.92 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.31 0.495 0.37 0.735 ;
        RECT 0.26 0.6 0.37 0.735 ;
        RECT 0.31 0.495 1.3 0.555 ;
        RECT 1.24 0.495 1.3 0.735 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END NAND3X2

MACRO ADDFHX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.745 0.415 4.805 0.555 ;
        RECT 4.745 1 4.805 1.39 ;
        RECT 4.745 0.495 5.285 0.555 ;
        RECT 5.155 1 5.215 1.39 ;
        RECT 5.165 0.415 5.225 0.555 ;
        RECT 5.225 0.495 5.285 1.06 ;
        RECT 4.745 1 5.285 1.06 ;
        RECT 5.225 0.6 5.34 0.73 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.28 0.6 0.34 0.98 ;
        RECT 0.34 0.52 0.4 0.66 ;
        RECT 0.34 0.92 0.4 1.295 ;
        RECT 0.28 0.92 0.82 0.98 ;
        RECT 0.76 0.52 0.82 0.66 ;
        RECT 0.26 0.6 0.82 0.66 ;
        RECT 0.76 0.92 0.82 1.295 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 0.79 2.525 0.85 ;
        RECT 2.26 0.79 2.525 0.94 ;
        RECT 2.26 0.88 3.235 0.94 ;
        RECT 3.175 0.82 4.325 0.88 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.54 0.63 1.6 0.75 ;
        RECT 1.54 0.63 2.685 0.69 ;
        RECT 2.625 0.63 2.685 0.78 ;
        RECT 2.625 0.72 3.075 0.78 ;
        RECT 3.015 0.66 4.485 0.72 ;
        RECT 4.235 0.625 4.485 0.72 ;
        RECT 4.425 0.625 4.485 0.745 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.435 2.365 0.53 ;
        RECT 2.235 0.47 2.825 0.53 ;
        RECT 2.795 0.5 2.915 0.62 ;
        RECT 2.765 0.5 4.015 0.56 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END ADDFHX4

MACRO NAND3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X4 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.415 1.015 0.475 1.405 ;
        RECT 0.825 1.125 0.885 1.405 ;
        RECT 1.235 1.125 1.295 1.405 ;
        RECT 1.645 1.125 1.705 1.405 ;
        RECT 2.055 1.125 2.115 1.405 ;
        RECT 0.415 1.125 2.525 1.185 ;
        RECT 2.465 1.04 2.525 1.405 ;
        RECT 0.895 0.405 2.74 0.465 ;
        RECT 2.66 0.98 2.74 1.11 ;
        RECT 2.68 0.405 2.74 1.11 ;
        RECT 2.465 1.05 2.74 1.11 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.815 0.365 0.895 ;
        RECT 0.305 0.855 0.7 0.915 ;
        RECT 0.64 0.855 0.7 1.025 ;
        RECT 1.475 0.885 1.595 1.025 ;
        RECT 2.305 0.88 2.365 1.025 ;
        RECT 0.64 0.965 2.365 1.025 ;
        RECT 2.495 0.82 2.555 0.94 ;
        RECT 2.305 0.88 2.555 0.94 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.515 0.695 0.86 0.755 ;
        RECT 0.8 0.695 0.86 0.865 ;
        RECT 1.265 0.725 1.325 0.865 ;
        RECT 0.8 0.805 1.325 0.865 ;
        RECT 1.265 0.725 1.755 0.785 ;
        RECT 1.695 0.725 1.755 0.865 ;
        RECT 2.145 0.685 2.205 0.865 ;
        RECT 1.695 0.805 2.205 0.865 ;
        RECT 2.26 0.6 2.34 0.745 ;
        RECT 2.26 0.625 2.395 0.745 ;
        RECT 2.145 0.685 2.395 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.565 1.165 0.705 ;
        RECT 0.96 0.645 1.165 0.705 ;
        RECT 1.035 0.565 1.915 0.625 ;
        RECT 1.855 0.565 1.915 0.705 ;
        RECT 1.855 0.645 1.985 0.705 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END NAND3X4

MACRO NOR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X8 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 0.995 0.715 1.385 ;
        RECT 1.3 0.995 1.36 1.385 ;
        RECT 2.195 0.995 2.255 1.385 ;
        RECT 0.655 0.995 3.14 1.055 ;
        RECT 2.915 0.96 2.975 1.385 ;
        RECT 0.32 0.49 3.14 0.55 ;
        RECT 3.08 0.49 3.14 1.11 ;
        RECT 2.915 0.96 3.14 1.11 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.69 0.81 0.91 0.87 ;
        RECT 1.41 0.81 1.53 0.895 ;
        RECT 2.025 0.81 2.145 0.895 ;
        RECT 2.635 0.815 2.93 0.86 ;
        RECT 0.85 0.835 2.765 0.895 ;
        RECT 2.705 0.8 2.93 0.86 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.78 0.54 0.84 ;
        RECT 0.48 0.65 0.54 0.92 ;
        RECT 0.46 0.78 0.54 0.92 ;
        RECT 1.01 0.65 1.13 0.735 ;
        RECT 1.805 0.65 1.925 0.735 ;
        RECT 0.48 0.65 2.305 0.71 ;
        RECT 2.245 0.675 2.565 0.735 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END NOR2X8

MACRO AOI32XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.88 0.425 0.94 1.11 ;
        RECT 0.86 0.98 0.94 1.11 ;
        RECT 0.86 1.05 1.26 1.11 ;
        RECT 1.2 1.05 1.26 1.245 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.48 0.48 0.56 0.89 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.23 1.14 0.73 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.22 0.74 0.35 ;
        RECT 0.665 0.27 0.745 0.715 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.72 1.34 0.92 ;
        RECT 1.26 0.84 1.44 0.92 ;
        RECT 1.36 0.84 1.44 1.12 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.62 0.34 1.12 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END AOI32XL

MACRO OAI22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.85 0.995 0.91 1.345 ;
        RECT 1.535 0.995 1.595 1.345 ;
        RECT 1.915 0.495 1.975 1.155 ;
        RECT 2.035 1.095 2.165 1.275 ;
        RECT 2.205 0.445 2.325 0.555 ;
        RECT 2.405 1.095 2.465 1.215 ;
        RECT 2.615 0.445 2.735 0.555 ;
        RECT 0.85 1.095 3.085 1.155 ;
        RECT 3.025 0.975 3.085 1.345 ;
        RECT 3.025 0.445 3.145 0.555 ;
        RECT 1.915 0.495 3.48 0.555 ;
        RECT 3.42 0.445 3.555 0.505 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.745 0.815 1.495 0.895 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.44 0.815 2.765 0.895 ;
        RECT 2.44 0.815 3.18 0.875 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.625 1.365 0.705 ;
        RECT 0.18 0.645 1.815 0.705 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.655 2.34 0.92 ;
        RECT 2.075 0.655 3.595 0.715 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END OAI22X4

MACRO OR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.87 0.395 0.94 1.085 ;
        RECT 0.86 0.79 0.94 1.085 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.53 0.59 0.61 0.91 ;
        RECT 0.53 0.79 0.74 0.91 ;
        RECT 0.66 0.79 0.74 0.96 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 0.96 ;
        RECT 0.19 0.59 0.27 0.87 ;
        RECT 0.06 0.79 0.27 0.87 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END OR2XL

MACRO SDFFSRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX4 0 0 ;
  SIZE 8.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 1.005 3.165 1.085 ;
        RECT 2.89 1.005 3.34 1.065 ;
        RECT 3.28 1.005 3.34 1.405 ;
        RECT 4.08 1.225 4.14 1.405 ;
        RECT 3.28 1.345 4.14 1.405 ;
        RECT 4.08 1.225 4.52 1.285 ;
        RECT 4.46 1.28 5.135 1.34 ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.46 0.625 8.4 0.705 ;
        RECT 8.32 0.625 8.4 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.835 0.805 8.135 0.965 ;
        RECT 7.715 0.835 8.135 0.965 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.86 0.625 6.94 1.085 ;
        RECT 6.86 0.865 6.98 1.085 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.435 0.815 6.76 0.895 ;
        RECT 6.68 0.815 6.76 1.07 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.75 1.74 1.25 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.54 0.495 1.29 ;
        RECT 0.435 0.625 0.565 0.705 ;
        RECT 0.435 0.645 0.86 0.705 ;
        RECT 0.8 0.585 0.86 0.96 ;
        RECT 0.845 0.525 0.905 0.645 ;
        RECT 0.845 0.9 0.905 1.29 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.6 0.06 ;
    END
  END VSS
END SDFFSRHQX4

MACRO TBUFX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX20 0 0 ;
  SIZE 10 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 0.475 5.945 0.66 ;
        RECT 5.885 0.6 6.14 0.66 ;
        RECT 5.975 1.05 6.035 1.415 ;
        RECT 6.02 0.6 6.08 1.11 ;
        RECT 6.02 0.6 6.14 0.73 ;
        RECT 6.295 0.475 6.355 0.615 ;
        RECT 6.385 0.555 6.445 1.415 ;
        RECT 6.705 0.475 6.765 0.615 ;
        RECT 6.295 0.555 6.765 0.615 ;
        RECT 6.795 1.025 6.855 1.415 ;
        RECT 7.115 0.475 7.175 0.615 ;
        RECT 7.205 0.555 7.265 1.415 ;
        RECT 7.525 0.475 7.585 0.615 ;
        RECT 7.115 0.555 7.585 0.615 ;
        RECT 7.615 1.025 7.675 1.415 ;
        RECT 7.935 0.475 7.995 0.615 ;
        RECT 8.025 1.025 8.085 1.415 ;
        RECT 7.935 0.555 8.405 0.615 ;
        RECT 8.345 0.475 8.405 1.085 ;
        RECT 8.435 1.025 8.495 1.415 ;
        RECT 8.755 0.475 8.815 0.615 ;
        RECT 8.845 1.025 8.905 1.415 ;
        RECT 9.165 0.475 9.225 0.615 ;
        RECT 9.255 1.025 9.315 1.415 ;
        RECT 9.575 0.475 9.68 0.615 ;
        RECT 8.755 0.555 9.68 0.615 ;
        RECT 6.02 1.025 9.725 1.085 ;
        RECT 9.62 0.475 9.68 1.085 ;
        RECT 9.665 1.025 9.725 1.415 ;
    END
  END Y
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.73 1.5 0.875 ;
        RECT 1.635 0.815 1.765 0.895 ;
        RECT 2 0.73 2.06 0.875 ;
        RECT 1.44 0.815 2.06 0.875 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.035 0.625 0.28 0.705 ;
        RECT 0.28 0.3 0.34 0.685 ;
        RECT 0.28 0.3 0.755 0.36 ;
        RECT 0.695 0.3 0.755 0.64 ;
        RECT 0.78 0.58 0.84 0.72 ;
        RECT 0.94 0.58 1 0.72 ;
        RECT 1.015 0.3 1.075 0.64 ;
        RECT 0.695 0.58 1.075 0.64 ;
        RECT 1.015 0.3 1.665 0.36 ;
        RECT 1.605 0.3 1.665 0.615 ;
        RECT 1.71 0.555 1.77 0.715 ;
        RECT 1.925 0.3 1.985 0.615 ;
        RECT 1.605 0.555 1.985 0.615 ;
        RECT 1.925 0.3 2.38 0.36 ;
        RECT 2.32 0.3 2.38 0.615 ;
        RECT 2.415 0.555 2.475 0.755 ;
        RECT 2.64 0.345 2.7 0.615 ;
        RECT 2.32 0.555 2.7 0.615 ;
        RECT 2.64 0.345 3.08 0.405 ;
        RECT 3.02 0.345 3.08 0.615 ;
        RECT 3.055 0.555 3.115 0.745 ;
        RECT 3.055 0.685 5.555 0.745 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 10 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 10 0.06 ;
    END
  END VSS
END TBUFX20

MACRO INVX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX16 0 0 ;
  SIZE 3.20 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.92 0.705 3 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.72 0.15 0.87 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.20 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.20 0.06 ;
    END
  END VSS
END INVX16

MACRO ADDHX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX4 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.08 0.815 3.14 1.25 ;
        RECT 3.28 0.57 3.34 0.92 ;
        RECT 3.26 0.79 3.34 0.92 ;
        RECT 3.08 0.815 3.695 0.875 ;
        RECT 3.07 0.57 3.66 0.63 ;
        RECT 3.635 0.815 3.695 1.02 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 0.52 0.86 0.64 ;
        RECT 1.26 0.58 1.34 1.01 ;
        RECT 0.91 0.95 1.34 1.01 ;
        RECT 1.28 0.58 1.34 1.13 ;
        RECT 1.44 0.51 1.5 0.64 ;
        RECT 0.8 0.58 1.5 0.64 ;
        RECT 1.28 1.07 1.5 1.13 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.2 0.92 ;
        RECT 0.14 0.76 0.2 1.2 ;
        RECT 0.14 1.14 0.88 1.2 ;
        RECT 0.82 1.14 0.88 1.29 ;
        RECT 0.82 1.23 1.98 1.29 ;
        RECT 1.92 0.78 1.98 1.435 ;
        RECT 1.905 0.78 2.025 0.84 ;
        RECT 1.92 1.375 2.745 1.435 ;
        RECT 2.685 1.35 3.3 1.41 ;
        RECT 3.24 1.12 3.3 1.41 ;
        RECT 3.88 0.74 3.94 1.18 ;
        RECT 3.24 1.12 3.94 1.18 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.54 0.8 ;
        RECT 0.64 0.36 0.7 0.66 ;
        RECT 0.46 0.6 0.7 0.66 ;
        RECT 0.64 0.36 1.34 0.42 ;
        RECT 1.28 0.35 1.66 0.41 ;
        RECT 1.6 0.35 1.66 0.68 ;
        RECT 1.6 0.62 1.855 0.68 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.2 0.06 ;
    END
  END VSS
END ADDHX4

MACRO SDFFSHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX8 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.54 0.335 1.345 ;
        RECT 0.685 0.54 0.745 1.345 ;
        RECT 0.275 0.6 1.155 0.66 ;
        RECT 1.06 0.6 1.155 0.73 ;
        RECT 1.095 0.54 1.155 1.345 ;
        RECT 1.505 0.93 1.565 1.05 ;
        RECT 1.62 0.54 1.68 0.99 ;
        RECT 1.095 0.93 1.68 0.99 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.045 0.73 7.92 0.79 ;
        RECT 7.86 0.79 7.94 0.92 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.32 0.945 7.76 1.085 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.235 0.7 6.365 0.905 ;
        RECT 6.235 0.81 6.61 0.89 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.015 0.755 6.135 0.835 ;
        RECT 6.035 0.755 6.135 1.085 ;
        RECT 6.035 1.005 6.265 1.085 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.435 1.005 2.565 1.085 ;
        RECT 2.505 0.93 2.565 1.35 ;
        RECT 2.505 0.93 2.575 1.05 ;
        RECT 3.515 1.22 3.575 1.35 ;
        RECT 2.505 1.29 3.575 1.35 ;
        RECT 3.775 0.95 3.835 1.28 ;
        RECT 3.515 1.22 3.835 1.28 ;
        RECT 3.775 0.95 3.94 1.01 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8 0.06 ;
    END
  END VSS
END SDFFSHQX8

MACRO DFFRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX2 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.53 0.34 1.305 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.815 1.715 1.115 ;
        RECT 1.485 1.025 1.715 1.115 ;
        RECT 1.635 0.815 1.765 0.895 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 0.74 0.765 1.085 ;
        RECT 0.6 1.005 0.835 1.085 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 0.515 4.175 0.705 ;
        RECT 4.095 0.515 4.175 0.885 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END DFFRHQX2

MACRO DFFNSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX4 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.79 6.34 0.92 ;
        RECT 6.48 0.86 6.54 1.33 ;
        RECT 6.595 0.505 6.655 0.92 ;
        RECT 6.26 0.86 6.95 0.92 ;
        RECT 6.89 0.86 6.95 1.33 ;
        RECT 6.595 0.505 7.185 0.565 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.635 1.005 5.695 1.33 ;
        RECT 5.635 1.005 5.765 1.085 ;
        RECT 5.715 0.505 5.775 1.065 ;
        RECT 5.635 1.005 6.13 1.065 ;
        RECT 6.07 1.005 6.13 1.33 ;
        RECT 5.655 0.505 6.245 0.565 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.885 0.63 2.965 0.895 ;
        RECT 2.805 0.815 2.965 0.895 ;
        RECT 2.885 0.63 3.12 0.71 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.625 2.365 0.745 ;
        RECT 2.235 0.665 2.695 0.745 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.76 0.54 1.26 ;
    END
  END D
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.76 0.34 1.26 ;
    END
  END CKN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.8 0.06 ;
    END
  END VSS
END DFFNSRX4

MACRO TLATNSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRX4 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.69 0.54 5.75 0.68 ;
        RECT 5.77 0.935 5.83 1.315 ;
        RECT 5.815 0.62 5.875 0.995 ;
        RECT 5.815 0.62 5.94 0.92 ;
        RECT 6.1 0.54 6.16 0.68 ;
        RECT 5.69 0.62 6.16 0.68 ;
        RECT 5.815 0.86 6.24 0.92 ;
        RECT 6.18 0.86 6.24 1.315 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.05 0.54 4.11 0.68 ;
        RECT 4.06 0.925 4.125 1.315 ;
        RECT 4.08 0.62 4.14 1.11 ;
        RECT 4.06 0.925 4.535 0.985 ;
        RECT 4.46 0.54 4.52 0.68 ;
        RECT 4.05 0.62 4.52 0.68 ;
        RECT 4.475 0.925 4.535 1.315 ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.085 0.795 3.205 0.855 ;
        RECT 3.145 0.795 3.205 0.935 ;
        RECT 3.145 0.875 3.695 0.935 ;
        RECT 3.635 0.785 3.765 0.895 ;
        RECT 3.635 0.785 3.79 0.845 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.695 1.74 1.195 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.815 0.89 0.875 ;
        RECT 0.83 0.215 0.89 0.895 ;
        RECT 0.635 0.815 0.89 0.895 ;
        RECT 0.83 0.215 1.525 0.275 ;
        RECT 1.465 0.215 1.525 0.36 ;
        RECT 1.465 0.3 2.935 0.36 ;
    END
  END RN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.7 0.34 1.2 ;
    END
  END GN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END TLATNSRX4

MACRO ADDFHX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.39 1.025 4.45 1.39 ;
        RECT 4.435 0.54 4.495 1.085 ;
        RECT 4.435 0.6 4.54 0.73 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.28 0.54 0.34 1.29 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.855 1.895 0.915 ;
        RECT 1.835 0.905 1.965 1.085 ;
        RECT 2.935 0.82 2.995 0.965 ;
        RECT 1.835 0.905 2.995 0.965 ;
        RECT 2.935 0.82 3.97 0.88 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.145 0.7 1.265 0.76 ;
        RECT 1.23 0.695 2.465 0.755 ;
        RECT 2.775 0.66 2.835 0.805 ;
        RECT 2.405 0.745 2.835 0.805 ;
        RECT 3.835 0.625 3.965 0.72 ;
        RECT 2.775 0.66 4.13 0.72 ;
        RECT 4.07 0.66 4.13 0.78 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.435 1.965 0.585 ;
        RECT 1.835 0.525 2.65 0.585 ;
        RECT 2.59 0.5 2.65 0.645 ;
        RECT 2.59 0.5 3.67 0.56 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END ADDFHX2

MACRO NOR4BBXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBXL 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.83 0.255 0.89 0.51 ;
        RECT 0.83 0.45 1.32 0.51 ;
        RECT 1.26 0.255 1.32 1.41 ;
        RECT 0.74 1.35 1.32 1.41 ;
        RECT 1.26 0.79 1.34 0.92 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.98 0.74 1.25 ;
        RECT 0.68 0.77 0.76 1.15 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.98 0.94 1.125 ;
        RECT 1.005 0.77 1.085 1.12 ;
        RECT 0.86 0.98 1.085 1.12 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.815 1.715 1.155 ;
        RECT 1.525 1.075 1.715 1.155 ;
        RECT 1.635 0.815 1.765 0.895 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.03 0.685 0.4 0.895 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END NOR4BBXL

MACRO NOR2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X6 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.435 0.335 0.555 ;
        RECT 0.58 1.025 0.64 1.335 ;
        RECT 0.685 0.435 0.745 0.555 ;
        RECT 1.095 0.435 1.155 0.555 ;
        RECT 1.225 1.025 1.285 1.335 ;
        RECT 1.505 0.435 1.565 0.555 ;
        RECT 1.915 0.435 1.975 0.555 ;
        RECT 1.915 1.025 1.975 1.335 ;
        RECT 0.275 0.495 2.38 0.555 ;
        RECT 2.26 0.98 2.34 1.11 ;
        RECT 2.32 0.495 2.38 1.085 ;
        RECT 0.58 1.025 2.38 1.085 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.615 0.815 0.835 0.875 ;
        RECT 1.155 0.815 1.275 0.915 ;
        RECT 0.775 0.855 1.885 0.915 ;
        RECT 1.835 0.815 2.06 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.215 0.79 0.34 0.85 ;
        RECT 0.28 0.655 0.34 0.92 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.935 0.655 1.055 0.755 ;
        RECT 1.55 0.655 1.67 0.755 ;
        RECT 0.28 0.655 2.22 0.715 ;
        RECT 2.16 0.655 2.22 0.88 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END NOR2X6

MACRO CLKBUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX8 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.225 0.505 0.285 0.625 ;
        RECT 0.225 0.93 0.285 1.375 ;
        RECT 0.26 0.565 0.32 0.99 ;
        RECT 0.26 0.565 0.34 0.73 ;
        RECT 0.635 0.93 0.695 1.375 ;
        RECT 0.605 0.55 0.725 0.625 ;
        RECT 1.045 0.93 1.105 1.375 ;
        RECT 1.015 0.55 1.135 0.625 ;
        RECT 0.225 0.93 1.515 0.99 ;
        RECT 0.225 0.565 1.455 0.625 ;
        RECT 1.455 0.93 1.515 1.375 ;
        RECT 1.41 0.55 1.545 0.61 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.06 0.6 2.14 1.1 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END CLKBUFX8

MACRO NOR2BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.035 0.49 0.095 1.055 ;
        RECT 0.035 0.815 0.165 0.895 ;
        RECT 0.275 0.43 0.335 0.55 ;
        RECT 0.535 0.995 0.595 1.36 ;
        RECT 0.685 0.43 0.745 0.55 ;
        RECT 0.035 0.995 1.215 1.055 ;
        RECT 1.095 0.43 1.155 0.55 ;
        RECT 1.155 0.995 1.215 1.36 ;
        RECT 1.505 0.43 1.565 0.55 ;
        RECT 0.035 0.49 1.565 0.55 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.815 1.25 0.895 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.98 1.54 1.11 ;
        RECT 1.69 0.81 1.77 1.06 ;
        RECT 1.46 0.98 1.77 1.06 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END NOR2BX4

MACRO TLATNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRX1 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.41 0.94 0.54 ;
        RECT 0.88 0.41 0.94 1.33 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.305 0.73 ;
        RECT 0.225 0.54 0.305 1.29 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.98 4.14 1.18 ;
        RECT 4.165 0.785 4.245 1.06 ;
        RECT 4.06 0.98 4.245 1.06 ;
    END
  END GN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 0.3 3.765 0.36 ;
        RECT 3.705 0.3 3.765 0.905 ;
        RECT 3.635 0.815 3.765 0.895 ;
        RECT 3.705 0.845 3.96 0.905 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.82 0.8 2.9 1.08 ;
        RECT 2.86 0.62 2.94 0.92 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.2 0.81 1.28 1.11 ;
        RECT 1.06 0.98 1.28 1.11 ;
        RECT 1.2 0.81 1.34 0.89 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END TLATNSRX1

MACRO AOI2BB1XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.45 0.14 0.92 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.06 0.86 0.315 0.92 ;
        RECT 0.255 0.86 0.315 1.385 ;
        RECT 0.315 0.285 0.375 0.51 ;
        RECT 0.08 0.45 0.375 0.51 ;
        RECT 0.315 0.285 0.45 0.345 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.98 0.54 1.26 ;
        RECT 0.47 0.77 0.55 1.06 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.77 0.73 1.26 ;
        RECT 0.65 0.98 0.74 1.26 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.45 1.14 0.95 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END AOI2BB1XL

MACRO NOR3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X8 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 1.09 1.06 1.21 ;
        RECT 2.25 1.09 2.31 1.21 ;
        RECT 3.765 1.09 3.825 1.21 ;
        RECT 1 1.09 4.97 1.15 ;
        RECT 4.91 0.9 4.97 1.345 ;
        RECT 5.025 0.275 5.085 1.085 ;
        RECT 4.91 0.9 5.085 1.085 ;
        RECT 0.34 0.275 5.16 0.335 ;
        RECT 4.91 1.005 5.165 1.085 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.31 0.73 0.37 0.895 ;
        RECT 0.235 0.815 0.37 0.895 ;
        RECT 0.235 0.835 0.575 0.895 ;
        RECT 0.515 0.835 0.575 0.99 ;
        RECT 1.625 0.77 1.745 0.83 ;
        RECT 1.685 0.77 1.745 0.99 ;
        RECT 2.83 0.77 2.89 0.99 ;
        RECT 2.83 0.77 2.95 0.83 ;
        RECT 4.19 0.77 4.25 0.99 ;
        RECT 0.515 0.93 4.25 0.99 ;
        RECT 4.19 0.77 4.31 0.83 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.675 0.735 0.735 ;
        RECT 0.675 0.675 0.735 0.83 ;
        RECT 1.205 0.62 1.265 0.83 ;
        RECT 0.675 0.77 1.265 0.83 ;
        RECT 1.205 0.62 1.325 0.68 ;
        RECT 1.91 0.61 1.97 0.73 ;
        RECT 1.265 0.61 2.185 0.67 ;
        RECT 2.125 0.61 2.185 0.83 ;
        RECT 2.56 0.62 2.62 0.83 ;
        RECT 2.125 0.77 2.62 0.83 ;
        RECT 2.56 0.62 2.68 0.68 ;
        RECT 2.62 0.61 3.295 0.67 ;
        RECT 3.235 0.62 3.595 0.68 ;
        RECT 3.535 0.62 3.595 0.83 ;
        RECT 3.915 0.62 3.975 0.83 ;
        RECT 3.535 0.77 3.975 0.83 ;
        RECT 3.915 0.62 4.09 0.68 ;
        RECT 4.03 0.61 4.47 0.67 ;
        RECT 4.41 0.625 4.765 0.685 ;
        RECT 4.635 0.625 4.765 0.705 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 0.435 1.07 0.67 ;
        RECT 2.345 0.435 2.405 0.67 ;
        RECT 2.285 0.61 2.405 0.67 ;
        RECT 3.695 0.435 3.755 0.67 ;
        RECT 3.695 0.61 3.815 0.67 ;
        RECT 0.835 0.435 4.925 0.495 ;
        RECT 4.865 0.435 4.925 0.725 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.2 0.06 ;
    END
  END VSS
END NOR3X8

MACRO ADDHX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX2 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.21 0.525 2.34 0.605 ;
        RECT 2.26 0.525 2.34 0.99 ;
        RECT 2.26 0.91 2.41 0.99 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.77 0.555 1.14 0.635 ;
        RECT 1.06 0.555 1.14 1.115 ;
        RECT 0.865 1.035 1.14 1.115 ;
    END
  END CO
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.615 0.895 0.765 1.085 ;
        RECT 0.705 0.895 0.765 1.275 ;
        RECT 0.705 1.215 0.91 1.275 ;
        RECT 0.85 1.215 0.91 1.34 ;
        RECT 0.85 1.28 1.36 1.34 ;
        RECT 1.3 1.28 1.36 1.4 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.365 0.32 0.83 ;
        RECT 0.26 0.6 0.34 0.83 ;
        RECT 1.46 0.365 1.52 0.96 ;
        RECT 1.71 0.23 1.83 0.425 ;
        RECT 0.26 0.365 2.785 0.425 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END ADDHX2

MACRO SDFFSHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX2 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.5 0.705 ;
        RECT 0.42 0.51 0.5 1.29 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.525 0.635 6.34 0.715 ;
        RECT 6.26 0.6 6.34 0.73 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.745 0.815 5.825 0.98 ;
        RECT 5.745 0.815 6.16 0.895 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.565 0.625 4.98 0.705 ;
        RECT 4.86 0.625 4.98 0.79 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.56 0.89 4.765 1.085 ;
        RECT 4.56 0.89 4.945 0.97 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.815 1.165 0.895 ;
        RECT 1.105 0.815 1.165 1.245 ;
        RECT 2.485 0.965 2.545 1.245 ;
        RECT 1.105 1.185 2.545 1.245 ;
        RECT 2.485 0.965 2.605 1.025 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END SDFFSHQX2

MACRO OAI32X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X4 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.905 1.155 0.965 1.275 ;
        RECT 2.155 1.155 2.215 1.275 ;
        RECT 2.435 1.155 2.565 1.275 ;
        RECT 2.855 0.685 2.915 1.215 ;
        RECT 3.065 0.485 3.125 0.745 ;
        RECT 2.855 0.685 3.125 0.745 ;
        RECT 3.065 0.485 3.185 0.595 ;
        RECT 3.25 1.155 3.31 1.275 ;
        RECT 3.475 0.485 3.595 0.595 ;
        RECT 0.905 1.155 3.93 1.215 ;
        RECT 3.87 1.155 3.93 1.275 ;
        RECT 3.885 0.485 4.005 0.595 ;
        RECT 3.065 0.535 4.34 0.595 ;
        RECT 4.28 0.485 4.415 0.545 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.815 0.38 0.895 ;
        RECT 0.32 0.815 0.38 1.055 ;
        RECT 1.425 0.885 1.545 1.055 ;
        RECT 2.695 0.855 2.755 1.055 ;
        RECT 0.32 0.995 2.755 1.055 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.015 0.845 3.075 1.055 ;
        RECT 3.595 0.885 3.715 1.055 ;
        RECT 4.115 0.855 4.175 1.055 ;
        RECT 3.015 0.995 4.175 1.055 ;
        RECT 4.26 0.79 4.34 0.92 ;
        RECT 4.115 0.855 4.34 0.92 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.815 0.765 0.895 ;
        RECT 1.265 0.725 1.325 0.875 ;
        RECT 0.48 0.815 1.325 0.875 ;
        RECT 1.265 0.725 1.86 0.785 ;
        RECT 1.8 0.725 1.86 0.895 ;
        RECT 1.8 0.835 2.585 0.895 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.295 0.725 3.895 0.785 ;
        RECT 3.835 0.775 4.005 0.895 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.625 1.165 0.705 ;
        RECT 0.915 0.645 1.165 0.705 ;
        RECT 1.105 0.565 2.075 0.625 ;
        RECT 2.015 0.565 2.075 0.735 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END OAI32X4

MACRO NAND4BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BXL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.3 0.14 0.54 ;
        RECT 0.08 0.3 0.14 1.12 ;
        RECT 0.215 0.24 0.275 0.36 ;
        RECT 0.06 0.3 0.275 0.36 ;
        RECT 0.34 1.06 0.46 1.215 ;
        RECT 0.08 1.06 0.62 1.12 ;
        RECT 0.56 1.06 0.62 1.215 ;
        RECT 0.56 1.155 0.86 1.215 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.775 1.115 1.225 ;
        RECT 1.035 0.775 1.165 0.895 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.23 0.74 0.73 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.25 0.54 0.73 ;
        RECT 0.46 0.6 0.56 0.73 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.46 0.34 0.96 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END NAND4BXL

MACRO TLATNCAX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX16 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 0.54 0.725 1.07 ;
        RECT 1.045 0.57 1.105 1.07 ;
        RECT 1.045 0.57 1.165 0.63 ;
        RECT 1.455 0.57 1.515 1.07 ;
        RECT 1.455 0.57 1.575 0.63 ;
        RECT 1.865 0.57 1.93 1.07 ;
        RECT 1.865 0.57 1.985 0.63 ;
        RECT 2.26 0.57 2.32 1.07 ;
        RECT 2.26 0.79 2.34 1.07 ;
        RECT 2.26 0.57 2.395 0.63 ;
        RECT 2.715 0.525 2.775 1.07 ;
        RECT 2.715 0.585 3.125 0.645 ;
        RECT 0.58 1.01 3.16 1.07 ;
        RECT 3.08 0.57 3.215 0.63 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.66 0.67 6.78 1.01 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.33 0.65 0.41 0.97 ;
        RECT 0.46 0.6 0.54 0.73 ;
        RECT 0.33 0.65 0.54 0.73 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.2 0.06 ;
    END
  END VSS
END TLATNCAX16

MACRO FILL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL1 0 0 ;
  SIZE 0.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.2 0.06 ;
    END
  END VSS
END FILL1

MACRO DFFSHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.54 0.34 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.465 0.71 4.77 0.79 ;
        RECT 4.635 0.71 4.77 0.985 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.235 0.71 4.365 1.05 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.35 1.52 0.92 ;
        RECT 1.17 0.86 1.52 0.92 ;
        RECT 1.46 0.6 1.54 0.73 ;
        RECT 1.46 0.35 2.72 0.41 ;
        RECT 2.66 0.35 2.72 0.705 ;
        RECT 2.66 0.645 2.94 0.705 ;
        RECT 2.88 0.645 2.94 0.82 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END DFFSHQX2

MACRO TBUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX3 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.97 1.11 2.03 1.23 ;
        RECT 2.04 0.4 2.1 0.54 ;
        RECT 2.26 0.48 2.32 1.17 ;
        RECT 1.97 1.11 2.32 1.17 ;
        RECT 2.26 0.79 2.34 0.96 ;
        RECT 2.26 0.9 2.5 0.96 ;
        RECT 2.44 0.9 2.5 1.29 ;
        RECT 2.45 0.4 2.51 0.54 ;
        RECT 2.04 0.48 2.51 0.54 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.83 0.965 0.89 ;
        RECT 0.835 0.27 0.895 0.895 ;
        RECT 0.835 0.815 0.965 0.895 ;
        RECT 0.835 0.27 1.735 0.33 ;
        RECT 1.675 0.27 1.735 0.69 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.77 ;
        RECT 0.26 0.65 0.735 0.73 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END TBUFX3

MACRO NOR2BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.48 0.14 0.92 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.49 0.46 0.61 0.54 ;
        RECT 0.06 0.86 0.76 0.92 ;
        RECT 0.7 0.86 0.76 1.36 ;
        RECT 0.08 0.48 0.98 0.54 ;
        RECT 0.93 0.46 1.05 0.52 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.98 1.14 1.14 ;
        RECT 1.22 0.8 1.3 1.06 ;
        RECT 1.06 0.98 1.3 1.06 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.8 0.94 1.3 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END NOR2BX2

MACRO AOI21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X4 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.785 0.445 0.905 0.505 ;
        RECT 1.405 0.445 1.525 0.525 ;
        RECT 1.89 0.465 1.95 0.895 ;
        RECT 1.95 0.405 2.01 0.525 ;
        RECT 1.89 0.815 2.165 0.895 ;
        RECT 2.06 0.815 2.165 1.075 ;
        RECT 0.855 0.465 2.395 0.525 ;
        RECT 2.345 0.445 2.465 0.505 ;
        RECT 2.06 0.955 2.53 1.015 ;
        RECT 2.47 0.955 2.53 1.075 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 0.815 1.45 0.895 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.54 0.655 1.74 0.715 ;
        RECT 1.66 0.655 1.74 0.92 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.625 2.365 0.715 ;
        RECT 2.05 0.635 2.54 0.715 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END AOI21X4

MACRO OR2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X6 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.225 0.96 1.285 1.43 ;
        RECT 1.3 0.35 1.36 0.66 ;
        RECT 1.635 0.96 1.695 1.43 ;
        RECT 1.71 0.35 1.77 0.66 ;
        RECT 1.86 0.6 1.92 1.02 ;
        RECT 1.86 0.6 1.94 0.73 ;
        RECT 1.225 0.96 2.105 1.02 ;
        RECT 2.045 0.96 2.105 1.43 ;
        RECT 2.12 0.35 2.18 0.66 ;
        RECT 1.3 0.6 2.18 0.66 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.91 0.54 1.3 ;
        RECT 0.46 0.91 0.665 0.99 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.77 0.34 0.92 ;
        RECT 0.26 0.77 0.36 0.85 ;
        RECT 0.28 0.73 0.965 0.81 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END OR2X6

MACRO OAI22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 1.025 0.7 1.355 ;
        RECT 0.935 0.625 0.995 1.085 ;
        RECT 0.835 1.005 0.995 1.085 ;
        RECT 1.1 0.445 1.16 0.685 ;
        RECT 0.935 0.625 1.16 0.685 ;
        RECT 1.1 0.445 1.245 0.555 ;
        RECT 0.64 1.025 1.465 1.085 ;
        RECT 1.405 1.025 1.465 1.355 ;
        RECT 1.1 0.495 1.58 0.555 ;
        RECT 1.52 0.445 1.655 0.505 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.805 0.34 1.11 ;
        RECT 0.26 0.805 0.655 0.885 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.835 1.74 0.915 ;
        RECT 1.66 0.835 1.74 1.115 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.2 0.625 0.835 0.705 ;
        RECT 0.755 0.625 0.835 0.745 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.095 0.785 1.34 0.865 ;
        RECT 1.26 0.655 1.34 0.92 ;
        RECT 1.26 0.655 1.73 0.735 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END OAI22X2

MACRO TBUFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX1 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.735 0.435 1.965 0.555 ;
        RECT 1.905 0.435 1.965 1.3 ;
        RECT 1.87 0.91 1.965 1.3 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.005 0.765 1.085 ;
        RECT 0.72 0.31 0.78 0.725 ;
        RECT 0.72 0.665 0.88 0.725 ;
        RECT 0.82 0.665 0.88 1.065 ;
        RECT 0.43 1.005 0.88 1.065 ;
        RECT 0.72 0.31 1.29 0.37 ;
        RECT 1.23 0.285 1.43 0.345 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 0.825 0.33 0.945 ;
        RECT 0.46 0.6 0.54 0.905 ;
        RECT 0.25 0.825 0.72 0.905 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END TBUFX1

MACRO SDFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX4 0 0 ;
  SIZE 7 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.67 0.49 5.74 1.29 ;
        RECT 5.66 0.79 5.74 1.29 ;
        RECT 5.66 0.9 6.15 0.96 ;
        RECT 6.09 0.9 6.15 1.29 ;
        RECT 5.67 0.49 6.26 0.55 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.86 0.79 4.92 1.29 ;
        RECT 4.88 0.49 4.94 0.96 ;
        RECT 4.86 0.9 5.33 0.96 ;
        RECT 4.73 0.49 5.32 0.55 ;
        RECT 5.27 0.9 5.33 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.64 1.765 0.72 ;
        RECT 1.635 0.64 1.765 0.895 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.38 1.34 0.88 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.98 0.54 1.17 ;
        RECT 0.58 0.79 0.66 1.11 ;
        RECT 0.46 0.98 0.66 1.11 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.395 0.57 0.475 0.69 ;
        RECT 0.26 0.6 0.84 0.69 ;
        RECT 0.76 0.6 0.84 0.96 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7 0.06 ;
    END
  END VSS
END SDFFX4

MACRO INVX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX12 0 0 ;
  SIZE 2.40 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 0.705 2.18 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.72 0.15 0.87 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.40 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.40 0.06 ;
    END
  END VSS
END INVX12

MACRO DFFRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX8 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.435 0.635 6.565 1.085 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.745 0.345 1.805 0.795 ;
        RECT 1.66 0.6 1.805 0.795 ;
        RECT 1.745 0.345 2.445 0.405 ;
        RECT 2.385 0.345 2.445 0.81 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.83 0.47 5.965 0.705 ;
        RECT 5.83 0.47 6.175 0.615 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.54 0.13 1.345 ;
        RECT 0.06 0.54 0.14 0.73 ;
        RECT 0.48 0.67 0.54 1.345 ;
        RECT 0.49 0.54 0.55 0.73 ;
        RECT 0.06 0.67 0.96 0.73 ;
        RECT 0.89 0.67 0.95 1.345 ;
        RECT 0.9 0.54 0.96 0.8 ;
        RECT 0.89 0.74 1.315 0.8 ;
        RECT 1.255 0.57 1.315 0.96 ;
        RECT 1.3 0.9 1.36 1.345 ;
        RECT 1.255 0.57 1.4 0.63 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END DFFRHQX8

MACRO NOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.435 0.495 0.555 ;
        RECT 0.74 0.995 0.8 1.345 ;
        RECT 0.845 0.435 0.905 0.555 ;
        RECT 1.255 0.435 1.315 0.555 ;
        RECT 1.405 0.995 1.465 1.345 ;
        RECT 1.665 0.435 1.725 0.555 ;
        RECT 0.435 0.495 1.965 0.555 ;
        RECT 1.835 0.815 1.965 0.895 ;
        RECT 1.905 0.495 1.965 1.055 ;
        RECT 0.74 0.995 1.965 1.055 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 0.815 1.42 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.655 0.54 0.92 ;
        RECT 0.365 0.655 1.795 0.715 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END NOR2X4

MACRO OR3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X8 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.905 1.695 1.345 ;
        RECT 1.705 0.57 1.825 0.63 ;
        RECT 2.045 0.905 2.105 1.345 ;
        RECT 2.115 0.57 2.235 0.645 ;
        RECT 2.455 0.905 2.515 1.345 ;
        RECT 2.555 0.525 2.615 0.645 ;
        RECT 2.66 0.585 2.72 0.965 ;
        RECT 2.66 0.585 2.74 0.73 ;
        RECT 1.635 0.905 2.925 0.965 ;
        RECT 2.865 0.905 2.925 1.345 ;
        RECT 1.78 0.585 2.98 0.645 ;
        RECT 2.935 0.57 3.055 0.63 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.825 0.74 1.11 ;
        RECT 0.66 0.825 0.955 0.905 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.53 0.665 1.195 0.725 ;
        RECT 1.06 0.665 1.14 0.92 ;
        RECT 1.06 0.665 1.195 0.785 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.52 0.34 0.73 ;
        RECT 0.295 0.505 1.36 0.565 ;
        RECT 1.3 0.505 1.36 0.755 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END OR3X8

MACRO BUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.365 0.73 ;
        RECT 0.305 0.555 0.365 0.925 ;
        RECT 0.35 0.495 0.41 0.615 ;
        RECT 0.35 0.865 0.41 1.32 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.76 0.765 1.085 ;
        RECT 0.51 1.005 0.765 1.085 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END BUFX2

MACRO NOR4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X8 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.455 0.38 0.515 ;
        RECT 0.67 0.455 0.79 0.53 ;
        RECT 1.08 0.455 1.2 0.53 ;
        RECT 1.49 0.455 1.61 0.53 ;
        RECT 1.95 0.455 2.07 0.53 ;
        RECT 2.36 0.455 2.48 0.53 ;
        RECT 2.77 0.455 2.89 0.53 ;
        RECT 3.18 0.455 3.3 0.53 ;
        RECT 3.59 0.455 3.71 0.53 ;
        RECT 4 0.455 4.12 0.53 ;
        RECT 4.41 0.455 4.53 0.53 ;
        RECT 4.645 0.995 4.705 1.185 ;
        RECT 4.82 0.455 4.94 0.53 ;
        RECT 5.055 0.995 5.115 1.185 ;
        RECT 5.23 0.455 5.35 0.53 ;
        RECT 5.3 0.815 5.525 1.055 ;
        RECT 4.645 0.995 5.525 1.055 ;
        RECT 5.46 0.79 5.525 1.185 ;
        RECT 5.3 0.815 5.54 0.92 ;
        RECT 5.49 0.47 5.55 0.875 ;
        RECT 5.67 0.41 5.73 0.53 ;
        RECT 0.335 0.47 5.73 0.53 ;
        RECT 5.3 0.815 5.935 0.875 ;
        RECT 5.875 0.815 5.935 1.345 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.75 0.94 0.92 ;
        RECT 0.95 0.71 1.03 0.83 ;
        RECT 0.4 0.75 1.03 0.83 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 0.77 2.165 0.895 ;
        RECT 1.885 0.77 2.545 0.85 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.32 0.77 4.34 0.83 ;
        RECT 4.225 0.71 4.285 0.83 ;
        RECT 4.26 0.77 4.34 0.92 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.755 0.63 4.965 0.895 ;
        RECT 4.755 0.63 5.39 0.71 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.2 0.06 ;
    END
  END VSS
END NOR4X8

MACRO AOI21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.625 1.36 0.74 ;
        RECT 1.46 0.485 1.565 0.705 ;
        RECT 1.24 0.625 1.565 0.705 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.59 0.865 0.67 ;
        RECT 0.66 0.59 0.74 0.73 ;
        RECT 0.66 0.59 0.865 0.71 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.77 0.56 0.9 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.505 0.41 0.625 0.47 ;
        RECT 0.575 0.43 1.14 0.49 ;
        RECT 1.06 0.43 1.14 0.73 ;
        RECT 1.08 0.37 1.14 0.9 ;
        RECT 1.08 0.84 1.265 0.9 ;
        RECT 1.205 0.84 1.265 1.02 ;
    END
  END Y
END AOI21X2

MACRO DFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.075 0.57 4.14 1.405 ;
        RECT 4.06 0.79 4.14 1.405 ;
        RECT 4.06 1.015 4.145 1.405 ;
        RECT 4.06 1.015 4.555 1.075 ;
        RECT 4.495 1.015 4.555 1.405 ;
        RECT 4.075 0.57 4.665 0.63 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.6 3.34 0.73 ;
        RECT 3.265 0.6 3.325 1.405 ;
        RECT 3.28 0.44 3.34 1.075 ;
        RECT 3.265 1.015 3.735 1.075 ;
        RECT 3.135 0.44 3.725 0.5 ;
        RECT 3.675 1.015 3.735 1.405 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.525 0.94 1.025 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.565 0.14 0.965 ;
        RECT 0.06 0.565 0.24 0.73 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END DFFX4

MACRO CLKBUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX12 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.475 0.295 1.04 ;
        RECT 0.28 0.255 0.34 0.535 ;
        RECT 0.26 0.98 0.34 1.45 ;
        RECT 0.69 0.255 0.75 0.535 ;
        RECT 0.69 0.98 0.75 1.45 ;
        RECT 1.1 0.255 1.16 0.535 ;
        RECT 1.1 0.98 1.16 1.45 ;
        RECT 1.51 0.255 1.57 0.535 ;
        RECT 1.51 0.98 1.57 1.45 ;
        RECT 0.235 0.98 1.98 1.04 ;
        RECT 1.92 0.255 1.98 0.535 ;
        RECT 0.235 0.475 1.98 0.535 ;
        RECT 1.92 0.98 1.98 1.45 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.795 2.34 1.23 ;
        RECT 2.26 0.795 2.405 0.875 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END CLKBUFX12

MACRO NOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X2 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 0.47 0.36 0.61 ;
        RECT 0.505 0.89 0.565 1.41 ;
        RECT 0.71 0.47 0.77 0.61 ;
        RECT 0.3 0.55 1.12 0.61 ;
        RECT 1.06 0.55 1.12 0.95 ;
        RECT 1.06 0.79 1.14 0.95 ;
        RECT 0.505 0.89 1.14 0.95 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.89 0.34 1.325 ;
        RECT 0.26 0.89 0.405 0.97 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.71 0.14 0.92 ;
        RECT 0.06 0.71 0.84 0.79 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END NOR2X2

MACRO TIELO
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELO 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.16 0.14 0.66 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.6 0.06 ;
    END
  END VSS
END TIELO

MACRO SDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX1 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.2 0.73 ;
        RECT 0.14 0.54 0.2 1.475 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.935 0.645 3.995 0.945 ;
        RECT 4.635 0.625 4.77 0.705 ;
        RECT 3.935 0.645 4.77 0.705 ;
        RECT 4.71 0.625 4.77 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.265 0.805 4.565 1.04 ;
        RECT 4.265 0.805 4.61 0.895 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 0.545 3.54 0.73 ;
        RECT 3.46 0.65 3.675 0.73 ;
        RECT 3.595 0.65 3.675 0.91 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 1.255 ;
        RECT 0.485 0.78 0.565 1.035 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END SDFFHQX1

MACRO NOR3BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX4 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.06 0.41 0.315 0.47 ;
        RECT 0.255 0.375 0.315 1.185 ;
        RECT 0.925 1.125 0.985 1.375 ;
        RECT 0.255 1.125 2.235 1.185 ;
        RECT 2.175 1.125 2.235 1.375 ;
        RECT 0.255 0.375 2.895 0.435 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 0.865 ;
        RECT 1.505 0.695 1.565 0.865 ;
        RECT 0.66 0.805 1.565 0.865 ;
        RECT 1.505 0.695 2 0.755 ;
        RECT 1.94 0.695 2 0.865 ;
        RECT 2.59 0.685 2.65 0.865 ;
        RECT 1.94 0.805 2.65 0.865 ;
        RECT 2.59 0.685 2.715 0.745 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.815 0.535 3.1 0.705 ;
        RECT 3.02 0.535 3.1 0.79 ;
        RECT 3.02 0.71 3.14 0.79 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.625 1.165 0.705 ;
        RECT 1.345 0.535 1.405 0.705 ;
        RECT 1.035 0.645 1.405 0.705 ;
        RECT 1.345 0.535 2.225 0.595 ;
        RECT 2.165 0.535 2.225 0.705 ;
        RECT 2.165 0.645 2.285 0.705 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END NOR3BX4

MACRO INVX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX3 0 0 ;
  SIZE 0.80 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 0.72 0.745 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.62 0.175 0.845 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.80 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.80 0.06 ;
    END
  END VSS
END INVX3

MACRO CLKXOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X4 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.435 0.32 1.29 ;
        RECT 0.26 0.435 0.335 0.575 ;
        RECT 0.26 0.79 0.335 1.29 ;
        RECT 0.26 0.79 0.34 0.96 ;
        RECT 0.26 0.9 0.7 0.96 ;
        RECT 0.64 0.355 0.7 0.575 ;
        RECT 0.26 0.515 0.7 0.575 ;
        RECT 0.64 0.9 0.7 1.215 ;
        RECT 0.685 0.295 0.745 0.415 ;
        RECT 0.685 1.155 0.745 1.275 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.9 0.615 2.34 0.695 ;
        RECT 2.26 0.615 2.34 0.92 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.96 0.675 1.165 0.895 ;
        RECT 0.96 0.675 1.32 0.755 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END CLKXOR2X4

MACRO DFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX1 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.88 0.4 0.94 1.11 ;
        RECT 0.86 0.98 0.94 1.11 ;
        RECT 0.86 1.05 1.09 1.11 ;
        RECT 1.02 0.34 1.08 0.46 ;
        RECT 0.88 0.4 1.08 0.46 ;
        RECT 1.03 1.05 1.09 1.17 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.29 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.4 0.46 6.48 0.85 ;
        RECT 6.46 0.41 6.54 0.54 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.68 0.605 5.76 0.87 ;
        RECT 5.68 0.79 5.94 0.87 ;
        RECT 5.86 0.79 5.94 0.925 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.235 0.625 3.365 0.705 ;
        RECT 3.305 0.3 3.365 0.865 ;
        RECT 2.265 0.805 3.365 0.865 ;
        RECT 3.305 0.3 4.005 0.36 ;
        RECT 3.945 0.3 4.005 0.92 ;
        RECT 3.945 0.86 4.855 0.92 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.285 0.72 1.365 0.895 ;
        RECT 1.04 0.815 1.365 0.895 ;
        RECT 1.285 0.72 1.445 0.8 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END DFFSRX1

MACRO AO21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X4 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.02 0.37 1.08 0.51 ;
        RECT 1.225 0.85 1.285 1.4 ;
        RECT 1.43 0.37 1.49 0.51 ;
        RECT 1.02 0.45 1.72 0.51 ;
        RECT 1.225 0.85 1.72 0.91 ;
        RECT 1.635 1.01 1.695 1.4 ;
        RECT 1.66 0.45 1.72 1.065 ;
        RECT 1.66 0.6 1.94 0.66 ;
        RECT 1.86 0.6 1.94 0.73 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.59 0.34 1.09 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.61 0.56 1.09 ;
        RECT 0.46 0.79 0.56 1.09 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 0.61 0.76 1.09 ;
        RECT 0.66 0.79 0.76 1.09 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END AO21X4

MACRO SDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRX2 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.22 0.57 1.28 1.29 ;
        RECT 1.22 0.57 1.34 0.63 ;
        RECT 1.22 0.79 1.34 0.92 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.62 0.57 0.74 0.63 ;
        RECT 0.66 0.57 0.72 1.29 ;
        RECT 0.66 0.57 0.74 0.73 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.22 6.34 0.35 ;
        RECT 6.265 0.27 6.345 0.73 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.085 0.645 6.165 1.095 ;
        RECT 6.035 1.005 6.165 1.095 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.605 0.645 5.685 0.895 ;
        RECT 5.605 0.79 5.765 0.895 ;
        RECT 5.605 0.79 5.935 0.87 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.79 4.34 0.965 ;
        RECT 4.48 0.685 4.56 0.91 ;
        RECT 4.26 0.79 4.56 0.91 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.6 1.74 1.1 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END SDFFTRX2

MACRO SDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX2 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.86 0.6 4.96 0.73 ;
        RECT 4.9 0.57 4.96 1.355 ;
        RECT 4.87 0.57 4.99 0.63 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.4 0.57 4.52 0.63 ;
        RECT 4.46 0.57 4.52 1.355 ;
        RECT 4.46 0.6 4.54 0.73 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.46 4.14 0.96 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.18 0.84 1.26 1.21 ;
        RECT 1.26 0.79 1.34 0.92 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.995 0.74 1.075 ;
        RECT 0.66 0.995 0.74 1.3 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.815 0.34 0.935 ;
        RECT 0.235 0.815 0.74 0.895 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END SDFFX2

MACRO NOR3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X4 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.915 1.125 0.975 1.375 ;
        RECT 2.165 1.125 2.225 1.375 ;
        RECT 0.255 0.375 2.92 0.435 ;
        RECT 2.86 0.375 2.92 1.185 ;
        RECT 0.915 1.125 2.92 1.185 ;
        RECT 2.86 0.41 2.94 0.54 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.08 0.79 0.14 1.01 ;
        RECT 0.08 0.95 0.575 1.01 ;
        RECT 1.525 0.855 1.645 1.025 ;
        RECT 2.64 0.825 2.7 1.025 ;
        RECT 0.515 0.965 2.7 1.025 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.49 0.79 0.735 0.85 ;
        RECT 1.365 0.695 1.425 0.865 ;
        RECT 0.675 0.805 1.425 0.865 ;
        RECT 1.365 0.695 1.83 0.755 ;
        RECT 1.77 0.695 1.83 0.82 ;
        RECT 2.31 0.67 2.37 0.82 ;
        RECT 1.77 0.76 2.37 0.82 ;
        RECT 2.46 0.6 2.54 0.73 ;
        RECT 2.31 0.67 2.54 0.73 ;
        RECT 2.47 0.6 2.54 0.79 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 0.535 0.985 0.705 ;
        RECT 0.835 0.625 0.985 0.705 ;
        RECT 0.925 0.535 2.055 0.595 ;
        RECT 1.995 0.535 2.055 0.66 ;
        RECT 1.995 0.6 2.115 0.66 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END NOR3X4

MACRO AOI31X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.91 0.535 1.97 0.675 ;
        RECT 2.32 0.535 2.38 0.675 ;
        RECT 2.73 0.535 2.79 0.675 ;
        RECT 2.945 0.995 3.005 1.115 ;
        RECT 3.14 0.535 3.2 0.675 ;
        RECT 2.945 0.995 3.54 1.055 ;
        RECT 3.41 0.995 3.47 1.115 ;
        RECT 3.46 0.615 3.52 1.11 ;
        RECT 3.46 0.98 3.54 1.11 ;
        RECT 3.55 0.535 3.61 0.675 ;
        RECT 1.91 0.615 3.61 0.675 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.385 0.695 0.515 0.775 ;
        RECT 0.435 0.695 0.515 0.895 ;
        RECT 0.435 0.815 0.845 0.895 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.205 0.695 1.325 0.895 ;
        RECT 1.205 0.805 1.365 0.895 ;
        RECT 1.205 0.805 1.665 0.885 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 0.775 3.165 0.895 ;
        RECT 2.9 0.775 3.36 0.855 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 0.815 2.535 0.895 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END AOI31X4

MACRO OAI32X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X2 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.81 1.025 0.87 1.365 ;
        RECT 1.235 1.005 1.5 1.085 ;
        RECT 0.81 1.025 1.5 1.085 ;
        RECT 1.44 0.505 1.5 1.305 ;
        RECT 1.73 0.455 1.85 0.565 ;
        RECT 1.44 1.245 1.925 1.305 ;
        RECT 1.865 1.245 1.925 1.365 ;
        RECT 1.44 0.505 2.185 0.565 ;
        RECT 2.125 0.455 2.26 0.515 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.845 0.54 1.125 ;
        RECT 0.46 0.845 0.76 0.925 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.665 1.16 0.745 ;
        RECT 0.86 0.665 0.94 0.92 ;
        RECT 0.86 0.665 1.16 0.785 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.825 1.94 1.145 ;
        RECT 1.84 0.825 2.1 0.905 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.505 0.295 0.73 ;
        RECT 0.235 0.505 1.34 0.565 ;
        RECT 1.26 0.505 1.34 0.73 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.665 1.74 0.92 ;
        RECT 1.6 0.665 2.3 0.725 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END OAI32X2

MACRO CLKXOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.085 0.52 0.145 0.73 ;
        RECT 0.06 0.6 0.145 0.73 ;
        RECT 0.14 0.67 0.2 1.29 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 0.835 1.035 0.895 ;
        RECT 1.235 0.815 1.365 0.895 ;
        RECT 0.975 0.815 1.535 0.875 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.73 0.54 1.23 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END CLKXOR2X1

MACRO NOR4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X6 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.33 0.35 0.39 0.64 ;
        RECT 0.74 0.35 0.8 0.64 ;
        RECT 1.15 0.35 1.21 0.64 ;
        RECT 1.615 0.35 1.675 0.64 ;
        RECT 2.025 0.35 2.085 0.64 ;
        RECT 2.545 0.35 2.605 0.64 ;
        RECT 2.955 0.35 3.015 0.64 ;
        RECT 3.365 0.35 3.425 0.64 ;
        RECT 3.59 0.92 3.65 1.21 ;
        RECT 3.87 0.35 3.93 0.64 ;
        RECT 3.59 1.09 4.125 1.15 ;
        RECT 4.065 0.92 4.125 1.21 ;
        RECT 0.33 0.58 4.34 0.64 ;
        RECT 4.26 0.58 4.32 0.98 ;
        RECT 4.28 0.35 4.34 0.73 ;
        RECT 4.065 0.92 4.535 0.98 ;
        RECT 4.475 0.9 4.535 1.37 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 0.75 0.74 0.83 ;
        RECT 0.66 0.74 0.74 0.92 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.76 1.575 0.895 ;
        RECT 1.39 0.76 1.835 0.84 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.59 0.74 3.14 0.82 ;
        RECT 3.06 0.74 3.14 0.92 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.835 0.74 3.965 0.895 ;
        RECT 3.7 0.74 4.125 0.82 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END NOR4X6

MACRO AOI222X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.76 0.38 0.82 0.52 ;
        RECT 1.375 1.2 1.435 1.32 ;
        RECT 1.45 0.41 1.72 0.52 ;
        RECT 0.76 0.46 1.72 0.52 ;
        RECT 1.66 0.41 1.72 1.26 ;
        RECT 1.66 0.98 1.74 1.26 ;
        RECT 1.375 1.2 1.74 1.26 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.62 0.76 0.92 ;
        RECT 0.68 0.62 0.76 1.1 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.62 1.54 1.1 ;
    END
  END C1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.49 0.34 0.99 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.755 0.94 0.92 ;
        RECT 0.88 0.86 1.095 1.1 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.195 0.79 1.275 1.225 ;
        RECT 1.195 0.79 1.34 0.92 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.545 0.715 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END AOI222X1

MACRO NAND4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X8 0 0 ;
  SIZE 6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.97 0.35 1.39 ;
        RECT 0.29 1.11 0.76 1.17 ;
        RECT 0.7 0.97 0.76 1.39 ;
        RECT 1.11 1.02 1.17 1.39 ;
        RECT 1.52 0.945 1.58 1.39 ;
        RECT 1.93 1.02 1.99 1.39 ;
        RECT 0.7 1.02 2.4 1.08 ;
        RECT 2.34 0.97 2.4 1.39 ;
        RECT 2.75 0.945 2.81 1.39 ;
        RECT 2.34 0.97 3.22 1.03 ;
        RECT 3.16 0.945 3.22 1.39 ;
        RECT 3.57 0.945 3.63 1.39 ;
        RECT 3.98 1.02 4.04 1.39 ;
        RECT 4.39 0.945 4.45 1.39 ;
        RECT 4.8 0.995 4.86 1.39 ;
        RECT 3.16 1.02 5.27 1.08 ;
        RECT 5.21 0.995 5.27 1.39 ;
        RECT 5.46 0.57 5.52 1.055 ;
        RECT 5.46 0.57 5.54 0.73 ;
        RECT 5.21 0.995 5.68 1.055 ;
        RECT 5.62 0.945 5.68 1.39 ;
        RECT 4.565 0.57 5.915 0.63 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 0.79 1.03 0.87 ;
        RECT 0.86 0.79 0.94 0.92 ;
        RECT 0.95 0.785 1.03 0.905 ;
        RECT 0.86 0.79 1.03 0.905 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.865 0.785 1.945 0.905 ;
        RECT 1.865 0.79 2.14 0.905 ;
        RECT 2.06 0.79 2.14 0.92 ;
        RECT 1.865 0.79 2.495 0.87 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.84 0.725 3.92 0.845 ;
        RECT 3.27 0.785 3.92 0.845 ;
        RECT 3.86 0.79 3.94 0.92 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.705 0.815 5.36 0.895 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6 0.06 ;
    END
  END VSS
END NAND4X8

MACRO SDFFSX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX4 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.87 0.97 6.93 1.09 ;
        RECT 6.915 0.655 6.975 1.03 ;
        RECT 6.915 0.655 7.565 0.715 ;
        RECT 7.505 0.655 7.565 0.85 ;
        RECT 7.505 0.79 7.74 0.85 ;
        RECT 7.66 0.79 7.74 0.92 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.235 0.815 7.405 1.055 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.365 0.815 6.61 0.895 ;
        RECT 6.53 0.815 6.61 1.15 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.94 1.005 6.365 1.085 ;
        RECT 6.285 0.995 6.43 1.075 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.295 3.12 0.875 ;
        RECT 2.645 0.815 3.12 0.875 ;
        RECT 3.06 0.6 3.14 0.73 ;
        RECT 3.06 0.295 4.14 0.355 ;
        RECT 4.08 0.295 4.14 0.42 ;
        RECT 4.08 0.36 4.435 0.42 ;
        RECT 4.375 0.36 4.435 0.67 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.6 1.565 0.73 ;
        RECT 1.505 0.54 1.565 1.405 ;
        RECT 1.46 0.67 1.975 0.73 ;
        RECT 1.915 0.54 1.975 1.405 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.54 0.335 1.29 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.26 0.86 0.745 0.92 ;
        RECT 0.685 0.54 0.745 1.29 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8 0.06 ;
    END
  END VSS
END SDFFSX4

MACRO DFFSHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX8 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.035 0.7 6.17 0.98 ;
        RECT 5.87 0.9 6.17 0.98 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.69 0.7 5.77 0.98 ;
        RECT 5.47 0.815 5.77 0.98 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.235 2.92 0.855 ;
        RECT 2.585 0.795 2.92 0.855 ;
        RECT 2.86 0.41 2.94 0.54 ;
        RECT 2.86 0.235 3.865 0.295 ;
        RECT 3.805 0.27 4.085 0.33 ;
        RECT 4.025 0.27 4.085 0.73 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.54 0.14 1.345 ;
        RECT 0.49 0.54 0.55 1.345 ;
        RECT 0.9 0.54 0.96 1.345 ;
        RECT 0.06 0.6 1.37 0.66 ;
        RECT 1.31 0.54 1.37 1.345 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.2 0.06 ;
    END
  END VSS
END DFFSHQX8

MACRO NOR4BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX4 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.88 0.475 0.94 0.615 ;
        RECT 1.29 0.475 1.35 0.615 ;
        RECT 1.635 0.555 1.695 1.085 ;
        RECT 1.7 0.475 1.76 0.615 ;
        RECT 1.635 0.995 1.765 1.085 ;
        RECT 2.11 0.475 2.17 0.615 ;
        RECT 2.52 0.475 2.58 0.615 ;
        RECT 2.93 0.475 2.99 0.615 ;
        RECT 3.34 0.475 3.4 0.615 ;
        RECT 3.545 0.995 3.605 1.135 ;
        RECT 3.75 0.475 3.81 0.615 ;
        RECT 0.88 0.555 3.81 0.615 ;
        RECT 1.635 0.995 4.015 1.055 ;
        RECT 3.955 0.995 4.015 1.135 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.06 0.65 0.285 0.73 ;
        RECT 0.205 0.65 0.285 0.955 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 0.815 2.295 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.595 0.715 2.675 0.895 ;
        RECT 2.595 0.815 3.15 0.895 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.415 0.715 3.495 0.895 ;
        RECT 3.415 0.815 3.97 0.895 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END NOR4BX4

MACRO CLKINVX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX3 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.415 0.54 0.475 0.68 ;
        RECT 0.415 0.9 0.475 1.29 ;
        RECT 0.46 0.62 0.54 0.96 ;
        RECT 0.415 0.9 0.885 0.96 ;
        RECT 0.825 0.54 0.885 0.68 ;
        RECT 0.415 0.62 0.885 0.68 ;
        RECT 0.825 0.9 0.885 1.29 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.62 0.315 0.945 ;
        RECT 0.06 0.725 0.315 0.945 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END CLKINVX3

MACRO SDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.47 0.81 4.53 0.93 ;
        RECT 4.5 0.655 4.56 0.87 ;
        RECT 5.035 0.625 5.165 0.715 ;
        RECT 4.5 0.655 5.165 0.715 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.82 0.815 5.06 0.985 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.79 3.94 0.92 ;
        RECT 3.86 0.84 4.21 0.92 ;
        RECT 4.13 0.75 4.21 0.93 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.69 0.34 1.19 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 1.075 ;
        RECT 0.525 0.54 0.585 0.85 ;
        RECT 1.005 0.54 1.065 1.075 ;
        RECT 0.46 1.015 1.065 1.075 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END SDFFHQX4

MACRO NOR3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X6 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.295 0.465 0.605 ;
        RECT 0.875 0.295 0.935 0.605 ;
        RECT 0.405 0.545 0.935 0.605 ;
        RECT 1.035 1.155 1.095 1.275 ;
        RECT 1.345 0.295 1.405 0.415 ;
        RECT 1.815 0.295 1.875 0.415 ;
        RECT 2.285 0.295 2.345 0.575 ;
        RECT 2.445 1.155 2.505 1.275 ;
        RECT 2.755 0.295 2.815 0.415 ;
        RECT 3.225 0.295 3.285 0.415 ;
        RECT 3.535 1.155 3.595 1.275 ;
        RECT 0.875 0.355 3.755 0.415 ;
        RECT 3.695 0.295 3.755 0.605 ;
        RECT 3.695 0.545 4.14 0.605 ;
        RECT 4.06 0.98 4.14 1.215 ;
        RECT 4.08 0.545 4.14 1.215 ;
        RECT 1.035 1.155 4.14 1.215 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.815 0.39 0.895 ;
        RECT 0.33 0.815 0.39 1.055 ;
        RECT 1.585 0.885 1.705 1.055 ;
        RECT 2.84 0.885 2.96 1.055 ;
        RECT 3.9 0.845 3.96 1.055 ;
        RECT 0.33 0.995 3.96 1.055 ;
        RECT 3.905 0.76 3.965 0.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.425 0.725 1.485 0.895 ;
        RECT 0.505 0.835 1.485 0.895 ;
        RECT 1.425 0.725 1.865 0.785 ;
        RECT 1.805 0.725 1.865 0.895 ;
        RECT 1.965 0.775 2.025 0.895 ;
        RECT 2.68 0.725 2.74 0.895 ;
        RECT 1.805 0.835 2.74 0.895 ;
        RECT 2.68 0.725 3.12 0.785 ;
        RECT 3.06 0.725 3.12 0.895 ;
        RECT 3.635 0.815 3.795 0.895 ;
        RECT 3.735 0.725 3.795 0.895 ;
        RECT 3.06 0.835 3.795 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.625 1.155 0.735 ;
        RECT 1.035 0.625 1.165 0.705 ;
        RECT 1.265 0.565 1.325 0.705 ;
        RECT 1.035 0.645 1.325 0.705 ;
        RECT 1.265 0.565 2.185 0.625 ;
        RECT 2.125 0.565 2.185 0.735 ;
        RECT 2.52 0.565 2.58 0.735 ;
        RECT 2.125 0.675 2.58 0.735 ;
        RECT 2.52 0.565 3.28 0.625 ;
        RECT 3.22 0.565 3.28 0.735 ;
        RECT 3.22 0.675 3.565 0.735 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.2 0.06 ;
    END
  END VSS
END NOR3X6

MACRO TLATNX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNX1 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.07 0.395 3.175 0.515 ;
        RECT 3.035 0.435 3.175 0.515 ;
        RECT 3.095 0.395 3.175 1.29 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.46 0.54 2.54 1.34 ;
    END
  END QN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 0.78 2.115 1.23 ;
        RECT 2.035 1.005 2.165 1.085 ;
    END
  END GN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.785 0.34 0.98 ;
        RECT 0.45 0.785 0.53 0.98 ;
        RECT 0.26 0.9 0.53 0.98 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END TLATNX1

MACRO AO21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.2 0.395 1.26 0.66 ;
        RECT 1.26 0.6 1.34 0.73 ;
        RECT 1.265 0.6 1.34 1.48 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.59 0.34 1.09 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.535 0.46 0.615 0.835 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 0.635 0.94 1.005 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END AO21X2

MACRO AOI31X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.335 1.54 0.395 ;
        RECT 1.46 0.6 1.54 0.73 ;
        RECT 1.48 0.275 1.54 1.005 ;
        RECT 1.505 0.945 1.565 1.065 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 0.815 1.055 0.935 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.655 0.54 0.92 ;
        RECT 0.375 0.655 1.055 0.715 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.215 0.495 0.275 0.695 ;
        RECT 0.215 0.495 1.215 0.555 ;
        RECT 1.155 0.495 1.215 0.73 ;
        RECT 1.155 0.6 1.34 0.73 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.495 1.94 0.995 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END AOI31X2

MACRO NOR3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.85 1.02 0.91 1.14 ;
        RECT 0.245 0.32 1.54 0.38 ;
        RECT 1.46 0.32 1.52 1.08 ;
        RECT 0.85 1.02 1.52 1.08 ;
        RECT 1.46 0.32 1.54 0.54 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.815 0.565 0.895 ;
        RECT 0.485 0.8 0.92 0.88 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.64 1.145 0.7 ;
        RECT 1.06 0.64 1.14 0.92 ;
        RECT 1.06 0.64 1.145 0.76 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.48 0.14 0.73 ;
        RECT 0.06 0.48 1.315 0.54 ;
        RECT 1.255 0.48 1.315 0.705 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END NOR3X2

MACRO NOR3BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.32 0.14 0.92 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.06 0.86 0.895 0.92 ;
        RECT 0.835 0.86 0.895 1.32 ;
        RECT 0.08 0.32 1.5 0.38 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.995 0.8 1.14 0.88 ;
        RECT 1.06 0.8 1.14 1.235 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 0.64 1.34 0.7 ;
        RECT 1.26 0.64 1.34 0.92 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 0.64 1.68 1.08 ;
        RECT 1.6 0.64 1.74 0.92 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END NOR3BX2

MACRO DFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRX1 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.41 0.94 0.54 ;
        RECT 0.88 0.41 0.94 0.95 ;
        RECT 0.9 0.89 0.96 1.34 ;
        RECT 0.86 0.41 0.975 0.53 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.29 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.365 4.54 0.865 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.79 4.14 0.92 ;
        RECT 4.06 0.79 4.32 0.87 ;
        RECT 4.24 0.735 4.32 1.005 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.98 1.14 1.11 ;
        RECT 1.26 0.78 1.34 1.06 ;
        RECT 1.06 0.98 1.34 1.06 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END DFFTRX1

MACRO TLATXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATXL 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.475 3.14 1.045 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.27 0.405 2.35 1.49 ;
        RECT 2.155 1.36 2.35 1.49 ;
    END
  END QN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.76 1.94 1.26 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.56 0.625 0.64 1.025 ;
        RECT 0.46 0.79 0.64 1.025 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END TLATXL

MACRO AO22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 0.47 1.365 0.53 ;
        RECT 1.45 0.915 1.51 1.305 ;
        RECT 1.685 0.47 1.805 0.55 ;
        RECT 1.315 0.49 1.92 0.55 ;
        RECT 1.45 0.915 1.92 0.975 ;
        RECT 1.86 0.49 1.92 1.305 ;
        RECT 1.86 0.6 1.94 0.73 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.815 1.12 0.895 ;
        RECT 1.035 0.815 1.12 1.085 ;
        RECT 1.035 1.005 1.31 1.085 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.52 0.34 1.02 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.52 0.74 1.02 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.52 0.56 1 ;
        RECT 0.46 0.79 0.56 1 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END AO22X4

MACRO NAND4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X6 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.92 0.49 1.37 ;
        RECT 0.84 0.9 0.9 1.37 ;
        RECT 0.43 1.09 1.31 1.15 ;
        RECT 1.25 0.9 1.31 1.37 ;
        RECT 1.8 1.02 1.86 1.37 ;
        RECT 2.285 0.9 2.345 1.37 ;
        RECT 2.695 0.92 2.755 1.37 ;
        RECT 1.25 1.02 3.225 1.08 ;
        RECT 3.165 0.95 3.225 1.37 ;
        RECT 3.165 0.95 3.635 1.01 ;
        RECT 3.575 0.9 3.635 1.37 ;
        RECT 3.825 0.52 3.885 0.64 ;
        RECT 3.575 1.09 4.125 1.15 ;
        RECT 4.065 0.92 4.125 1.37 ;
        RECT 3.825 0.58 4.32 0.64 ;
        RECT 4.26 0.52 4.32 1.08 ;
        RECT 4.26 0.79 4.34 0.92 ;
        RECT 4.065 1.02 4.535 1.08 ;
        RECT 4.475 0.9 4.535 1.37 ;
        RECT 4.68 0.35 4.74 0.66 ;
        RECT 4.26 0.6 4.74 0.66 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.385 0.74 0.74 0.82 ;
        RECT 0.66 0.74 0.74 0.965 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.74 1.74 0.92 ;
        RECT 1.66 0.77 2.06 0.85 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.735 0.74 2.915 0.82 ;
        RECT 2.86 0.77 2.94 0.92 ;
        RECT 3.015 0.73 3.095 0.85 ;
        RECT 2.835 0.77 3.095 0.85 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.735 0.815 3.965 0.895 ;
        RECT 3.86 0.74 4.16 0.82 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END NAND4X6

MACRO SDFFSX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX2 0 0 ;
  SIZE 6.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.6 1.145 0.73 ;
        RECT 1.065 0.54 1.145 1.29 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.28 0.54 0.34 1.29 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.89 0.645 5.95 1.085 ;
        RECT 5.83 1.025 5.95 1.085 ;
        RECT 6.105 0.585 6.165 0.705 ;
        RECT 5.89 0.645 6.365 0.705 ;
        RECT 6.105 0.625 6.505 0.685 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.435 0.815 6.61 1.055 ;
        RECT 6.27 0.975 6.61 1.055 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.46 0.55 5.54 0.765 ;
        RECT 5.265 0.55 5.63 0.63 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.045 0.635 5.165 1.085 ;
        RECT 5.035 1.005 5.165 1.085 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.315 2.295 0.895 ;
        RECT 2.235 0.815 2.365 0.895 ;
        RECT 1.855 0.835 2.365 0.895 ;
        RECT 2.235 0.315 3.065 0.375 ;
        RECT 3.005 0.315 3.065 0.55 ;
        RECT 3.385 0.33 3.445 0.55 ;
        RECT 3.005 0.49 3.445 0.55 ;
        RECT 3.385 0.33 3.505 0.39 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.8 0.06 ;
    END
  END VSS
END SDFFSX2

MACRO MX3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.37 0.705 ;
        RECT 0.31 0.46 0.37 0.95 ;
        RECT 0.355 0.4 0.415 0.52 ;
        RECT 0.355 0.89 0.415 1.48 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.405 1.025 2.485 1.155 ;
        RECT 2.86 0.98 2.94 1.155 ;
        RECT 2.405 1.075 2.94 1.155 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.395 0.74 2.74 0.82 ;
        RECT 2.66 0.74 2.74 0.975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.79 1.94 0.985 ;
        RECT 1.895 0.52 1.975 0.87 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.52 1.74 1.02 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.71 0.78 0.79 1.085 ;
        RECT 0.515 1.005 0.79 1.085 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END MX3X2

MACRO NOR4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.59 0.515 0.65 0.655 ;
        RECT 1 0.515 1.06 0.655 ;
        RECT 1.06 0.79 1.14 0.92 ;
        RECT 1.08 0.595 1.14 1.055 ;
        RECT 1.41 0.515 1.47 0.655 ;
        RECT 1.82 0.515 1.88 0.655 ;
        RECT 2.23 0.515 2.29 0.655 ;
        RECT 2.64 0.515 2.7 0.655 ;
        RECT 2.995 0.995 3.055 1.135 ;
        RECT 3.05 0.515 3.11 0.655 ;
        RECT 1.08 0.995 3.465 1.055 ;
        RECT 3.405 0.995 3.465 1.135 ;
        RECT 3.46 0.515 3.52 0.655 ;
        RECT 0.59 0.595 3.52 0.655 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.755 0.94 0.95 ;
        RECT 0.35 0.87 0.94 0.95 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.725 0.755 1.805 0.895 ;
        RECT 1.24 0.815 1.805 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.435 0.775 2.57 0.895 ;
        RECT 2.11 0.815 2.57 0.895 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.105 0.775 3.185 0.895 ;
        RECT 2.835 0.815 3.42 0.895 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END NOR4X4

MACRO OAI222XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 1.23 0.81 1.385 ;
        RECT 1.395 0.305 1.455 0.515 ;
        RECT 1.395 0.455 1.5 0.515 ;
        RECT 1.46 1.23 1.555 1.49 ;
        RECT 1.44 0.47 1.7 0.53 ;
        RECT 1.64 0.47 1.7 1.29 ;
        RECT 0.75 1.23 1.7 1.29 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.63 0.94 1.13 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.63 0.34 1.13 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.61 1.34 1.11 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.765 0.54 1.26 ;
        RECT 0.46 0.765 0.545 0.92 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.63 1.54 1.13 ;
    END
  END C1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.63 1.14 1.13 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OAI222XL

MACRO AOI222X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.76 0.475 0.88 0.535 ;
        RECT 1.38 0.475 1.5 0.555 ;
        RECT 1.835 0.815 1.965 0.895 ;
        RECT 1.905 0.495 1.965 1.055 ;
        RECT 2.345 0.475 2.465 0.555 ;
        RECT 3.21 0.475 3.33 0.555 ;
        RECT 3.855 0.995 3.915 1.135 ;
        RECT 3.98 0.475 4.1 0.555 ;
        RECT 4.265 0.995 4.325 1.135 ;
        RECT 0.83 0.495 4.56 0.555 ;
        RECT 4.51 0.475 4.72 0.535 ;
        RECT 4.675 0.995 4.735 1.135 ;
        RECT 1.905 0.995 5.145 1.055 ;
        RECT 5.085 0.995 5.145 1.135 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.465 0.815 3.2 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.815 1.425 0.895 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.055 0.815 4.795 0.895 ;
    END
  END C1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.655 2.295 0.895 ;
        RECT 2.235 0.815 2.365 0.895 ;
        RECT 2.11 0.655 3.61 0.715 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.835 0.625 4.965 0.715 ;
        RECT 3.745 0.655 5.15 0.715 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.625 0.565 0.715 ;
        RECT 0.42 0.655 1.735 0.715 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END AOI222X4

MACRO CLKINVX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX6 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.9 0.335 1.37 ;
        RECT 0.285 0.245 0.345 0.525 ;
        RECT 0.275 1.09 0.755 1.15 ;
        RECT 0.695 0.245 0.755 0.525 ;
        RECT 0.695 0.9 0.755 1.37 ;
        RECT 0.86 0.465 0.92 0.96 ;
        RECT 0.86 0.79 0.94 0.96 ;
        RECT 0.695 0.9 1.165 0.96 ;
        RECT 1.105 0.245 1.165 0.525 ;
        RECT 0.285 0.465 1.165 0.525 ;
        RECT 1.105 0.9 1.165 1.37 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.625 0.73 0.705 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END CLKINVX6

MACRO NOR4BBX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX2 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.4 1.38 0.46 ;
        RECT 1.33 0.45 2.72 0.48 ;
        RECT 1.715 0.36 1.775 0.51 ;
        RECT 1.26 0.42 1.775 0.46 ;
        RECT 2.125 0.37 2.185 0.51 ;
        RECT 2.535 0.37 2.595 0.51 ;
        RECT 1.715 0.45 2.72 0.51 ;
        RECT 2.635 0.805 2.695 1.145 ;
        RECT 2.66 0.45 2.72 0.865 ;
        RECT 2.66 0.6 2.74 0.73 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.225 0.65 2.365 0.895 ;
        RECT 2.225 0.65 2.56 0.73 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 0.61 2.125 0.925 ;
        RECT 1.86 0.755 2.125 0.925 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.515 0.805 0.595 1.085 ;
        RECT 0.295 1.005 0.595 1.085 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 0.625 0.375 0.905 ;
        RECT 0.295 0.625 0.595 0.705 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END NOR4BBX2

MACRO OR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 0.885 0.895 1.29 ;
        RECT 0.84 0.38 0.9 0.5 ;
        RECT 0.86 0.45 0.92 0.94 ;
        RECT 0.86 0.6 0.94 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.73 0.51 1.14 ;
        RECT 0.43 0.73 0.535 0.895 ;
        RECT 0.43 0.815 0.6 0.895 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.36 0.14 0.54 ;
        RECT 0.09 0.46 0.17 0.83 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END OR2X1

MACRO MX4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.185 0.6 4.245 0.72 ;
        RECT 4.9 0.6 4.96 0.75 ;
        RECT 4.185 0.6 5.14 0.66 ;
        RECT 5.06 0.6 5.14 0.73 ;
    END
  END S0
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.405 0.815 4.485 1 ;
        RECT 4.405 0.815 4.8 0.895 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.465 0.805 3.545 1.085 ;
        RECT 3.465 1.005 3.765 1.085 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.235 0.805 3.365 1.115 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.46 0.53 2.54 1.03 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 0.435 1.325 0.85 ;
        RECT 1.235 0.435 1.4 0.515 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.435 1.72 0.99 ;
        RECT 1.66 0.77 1.74 0.99 ;
        RECT 1.66 0.86 1.75 0.99 ;
        RECT 1.63 0.93 1.75 0.99 ;
        RECT 1.66 0.86 2.16 0.92 ;
        RECT 2.1 0.465 2.16 0.99 ;
        RECT 2.1 0.465 2.22 0.525 ;
        RECT 2.1 0.93 2.22 0.99 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END MX4X4

MACRO MDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX1 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.2 0.73 ;
        RECT 0.14 0.54 0.2 1.475 ;
    END
  END Q
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.935 0.645 3.995 0.945 ;
        RECT 4.635 0.625 4.77 0.705 ;
        RECT 3.935 0.645 4.77 0.705 ;
        RECT 4.71 0.625 4.77 0.745 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.265 0.805 4.565 1.04 ;
        RECT 4.265 0.805 4.61 0.895 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 0.545 3.54 0.73 ;
        RECT 3.46 0.65 3.675 0.73 ;
        RECT 3.595 0.65 3.675 0.91 ;
    END
  END D0
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 1.255 ;
        RECT 0.485 0.78 0.565 1.035 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END MDFFHQX1

MACRO NOR4BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX2 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.985 0.405 1.045 0.545 ;
        RECT 1.26 0.79 1.355 0.92 ;
        RECT 1.295 0.485 1.355 1.055 ;
        RECT 1.395 0.405 1.455 0.545 ;
        RECT 1.845 0.405 1.905 0.545 ;
        RECT 2.255 0.405 2.315 0.545 ;
        RECT 0.985 0.485 2.315 0.545 ;
        RECT 1.295 0.995 2.52 1.055 ;
        RECT 2.46 0.995 2.52 1.135 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.36 0.735 0.455 0.87 ;
        RECT 0.06 0.79 0.455 0.87 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 0.645 1.535 0.895 ;
        RECT 1.635 0.8 1.77 0.895 ;
        RECT 1.455 0.815 1.77 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.87 0.645 2.035 0.895 ;
        RECT 1.87 0.815 2.2 0.895 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.3 0.645 2.565 0.895 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END NOR4BX2

MACRO DFFSRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX4 0 0 ;
  SIZE 7.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 1.005 3.165 1.085 ;
        RECT 2.975 1.005 3.425 1.065 ;
        RECT 3.365 1.005 3.425 1.405 ;
        RECT 4.165 1.225 4.225 1.405 ;
        RECT 3.365 1.345 4.225 1.405 ;
        RECT 4.165 1.225 4.605 1.285 ;
        RECT 4.545 1.28 5.205 1.34 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.005 0.625 7.085 0.84 ;
        RECT 7.005 0.625 7.37 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.275 0.815 6.585 0.945 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.605 0.625 1.775 0.865 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.415 0.495 1.34 ;
        RECT 0.435 0.6 0.54 0.73 ;
        RECT 0.435 0.67 0.905 0.73 ;
        RECT 0.845 0.415 0.905 1.34 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.4 0.06 ;
    END
  END VSS
END DFFSRHQX4

MACRO NAND4BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX2 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.115 0.945 1.395 ;
        RECT 1.18 0.655 1.24 1.175 ;
        RECT 1.26 1.115 1.355 1.3 ;
        RECT 1.295 1.115 1.355 1.395 ;
        RECT 1.705 1.115 1.765 1.395 ;
        RECT 0.885 1.115 2.205 1.175 ;
        RECT 2.115 1.115 2.205 1.395 ;
        RECT 2.22 0.455 2.28 0.715 ;
        RECT 1.18 0.655 2.28 0.715 ;
        RECT 2.22 0.455 2.355 0.515 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.03 0.705 0.26 0.79 ;
        RECT 0.18 0.705 0.26 0.895 ;
        RECT 0.18 0.815 0.42 0.895 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.34 0.815 1.565 1.015 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.665 0.815 1.965 1.015 ;
        RECT 1.665 0.85 2.045 1.015 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.16 0.815 2.57 0.97 ;
        RECT 2.145 0.89 2.57 0.97 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END NAND4BX2

MACRO AOI2BB1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 0.465 0.235 1.255 ;
        RECT 0.235 1.195 0.365 1.275 ;
        RECT 0.405 0.385 0.465 0.525 ;
        RECT 0.61 1.195 0.67 1.475 ;
        RECT 0.815 0.385 0.875 0.525 ;
        RECT 0.175 1.195 1.29 1.255 ;
        RECT 1.225 0.385 1.285 0.525 ;
        RECT 1.23 1.195 1.29 1.475 ;
        RECT 1.635 0.385 1.695 0.525 ;
        RECT 0.175 0.465 1.695 0.525 ;
    END
  END Y
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.435 1.94 0.935 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.5 2.34 1 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.785 0.54 0.92 ;
        RECT 0.335 0.785 1.755 0.845 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END AOI2BB1X4

MACRO AO22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.415 1.52 1.11 ;
        RECT 1.465 0.98 1.54 1.48 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 0.655 1.105 1.12 ;
        RECT 1.025 0.955 1.14 1.12 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.63 0.16 1.11 ;
        RECT 0.06 0.955 0.16 1.11 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.605 0.765 0.705 ;
        RECT 0.685 0.605 0.765 1.055 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.26 0.815 0.535 0.895 ;
        RECT 0.455 0.815 0.535 1.07 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END AO22X2

MACRO NOR4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.445 0.395 0.505 ;
        RECT 0.715 0.445 0.835 0.525 ;
        RECT 1.155 0.445 1.275 0.525 ;
        RECT 1.595 0.445 1.715 0.525 ;
        RECT 0.345 0.465 1.94 0.525 ;
        RECT 1.86 1.17 1.94 1.345 ;
        RECT 1.88 0.465 1.94 1.345 ;
        RECT 1.01 1.285 1.94 1.345 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.82 0.32 1.185 ;
        RECT 1.66 0.98 1.74 1.185 ;
        RECT 1.68 0.82 1.74 1.185 ;
        RECT 0.26 1.125 1.74 1.185 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 0.835 0.54 0.895 ;
        RECT 0.46 0.79 0.54 0.92 ;
        RECT 0.48 0.79 0.54 1.025 ;
        RECT 1.435 0.845 1.495 1.025 ;
        RECT 0.48 0.965 1.495 1.025 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.275 0.625 1.335 0.865 ;
        RECT 0.64 0.805 1.335 0.865 ;
        RECT 1.275 0.625 1.565 0.705 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.625 1.14 0.705 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END NOR4X2

MACRO DFFQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX1 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.175 0.73 ;
        RECT 0.095 0.48 0.175 1.44 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.76 1.005 2.965 1.175 ;
        RECT 2.76 1.005 3.17 1.085 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.72 0.54 1.22 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END DFFQX1

MACRO MX2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.26 1.52 1.385 ;
        RECT 1.46 0.98 1.54 1.11 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 0.84 1.295 1.245 ;
        RECT 1.26 0.79 1.34 0.92 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.495 0.615 0.575 1.08 ;
        RECT 0.46 0.79 0.575 1.08 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.36 1.11 ;
        RECT 0.28 0.98 0.36 1.26 ;
        RECT 0.675 1.005 0.755 1.26 ;
        RECT 0.28 1.18 0.755 1.26 ;
        RECT 0.675 1.005 0.795 1.085 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END MX2XL

MACRO XOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.085 0.52 0.145 0.73 ;
        RECT 0.06 0.6 0.145 0.73 ;
        RECT 0.14 0.67 0.2 1.29 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 0.835 1.035 0.895 ;
        RECT 1.235 0.815 1.365 0.895 ;
        RECT 0.975 0.815 1.535 0.875 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.73 0.54 1.23 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END XOR2X1

MACRO NAND4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X4 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.975 0.335 1.365 ;
        RECT 0.695 0.975 0.755 1.365 ;
        RECT 1.08 0.655 1.14 1.11 ;
        RECT 1.06 0.995 1.19 1.11 ;
        RECT 0.275 0.975 1.14 1.035 ;
        RECT 1.13 0.995 1.19 1.365 ;
        RECT 1.54 0.995 1.6 1.365 ;
        RECT 1.985 0.995 2.045 1.365 ;
        RECT 2.395 0.995 2.455 1.365 ;
        RECT 2.745 0.525 2.805 0.715 ;
        RECT 1.08 0.655 2.805 0.715 ;
        RECT 2.97 0.995 3.03 1.365 ;
        RECT 3.205 0.445 3.265 0.585 ;
        RECT 1.06 0.995 3.44 1.055 ;
        RECT 3.38 0.995 3.44 1.365 ;
        RECT 3.635 0.445 3.695 0.585 ;
        RECT 2.745 0.525 3.695 0.585 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.625 0.73 0.705 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.815 1.74 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.835 0.815 2.965 0.895 ;
        RECT 2.905 0.685 2.965 0.895 ;
        RECT 2.095 0.835 2.965 0.895 ;
        RECT 2.905 0.685 3.025 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.465 0.685 3.545 0.895 ;
        RECT 3.105 0.815 3.545 0.895 ;
        RECT 3.465 0.685 3.585 0.765 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END NAND4X4

MACRO AOI2BB1X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.435 0.14 0.815 ;
        RECT 0.08 0.755 0.31 0.815 ;
        RECT 0.25 0.755 0.31 1.475 ;
        RECT 0.08 0.435 0.42 0.495 ;
        RECT 0.37 0.415 0.49 0.475 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.98 0.54 1.235 ;
        RECT 0.48 0.755 0.56 1.06 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.755 0.74 1.255 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.67 1.08 1.06 ;
        RECT 1.06 0.98 1.14 1.11 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END AOI2BB1X1

MACRO CLKINVX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX16 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.995 0.465 1.345 ;
        RECT 0.375 0.57 0.495 0.63 ;
        RECT 0.815 0.995 0.895 1.345 ;
        RECT 0.785 0.57 0.905 0.645 ;
        RECT 1.225 0.995 1.285 1.345 ;
        RECT 1.195 0.57 1.315 0.645 ;
        RECT 0.405 0.995 1.695 1.055 ;
        RECT 1.635 0.93 1.695 1.345 ;
        RECT 1.605 0.57 1.725 0.645 ;
        RECT 2.045 0.93 2.105 1.345 ;
        RECT 2.015 0.57 2.135 0.645 ;
        RECT 2.455 0.93 2.515 1.345 ;
        RECT 2.425 0.57 2.545 0.645 ;
        RECT 2.865 0.525 2.925 0.645 ;
        RECT 0.45 0.585 2.97 0.645 ;
        RECT 2.865 0.93 2.925 1.345 ;
        RECT 2.86 0.93 2.94 1.11 ;
        RECT 2.91 0.585 2.97 0.99 ;
        RECT 1.635 0.93 2.97 0.99 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.77 0.765 0.895 ;
        RECT 0.515 0.77 2.81 0.83 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END CLKINVX16

MACRO BUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX8 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.225 0.505 0.285 0.625 ;
        RECT 0.225 0.93 0.285 1.375 ;
        RECT 0.26 0.565 0.32 0.99 ;
        RECT 0.26 0.565 0.34 0.73 ;
        RECT 0.635 0.93 0.695 1.375 ;
        RECT 0.605 0.55 0.725 0.625 ;
        RECT 1.045 0.93 1.105 1.375 ;
        RECT 1.015 0.55 1.135 0.625 ;
        RECT 0.225 0.93 1.515 0.99 ;
        RECT 0.225 0.565 1.455 0.625 ;
        RECT 1.455 0.93 1.515 1.375 ;
        RECT 1.41 0.55 1.545 0.61 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.06 0.6 2.14 1.1 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END BUFX8

MACRO AND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.82 0.53 0.965 0.705 ;
        RECT 0.87 0.53 0.965 1.48 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.77 0.55 1.26 ;
        RECT 0.46 0.98 0.55 1.26 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.12 0.8 0.2 1.23 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END AND2X1

MACRO NAND4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X2 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.32 1.285 0.38 1.405 ;
        RECT 0.79 1.285 0.85 1.405 ;
        RECT 1.07 0.445 1.235 0.505 ;
        RECT 1.26 1.285 1.32 1.405 ;
        RECT 1.73 1.285 1.79 1.405 ;
        RECT 1.185 0.465 2.12 0.525 ;
        RECT 2.06 0.465 2.12 1.345 ;
        RECT 2.06 1.17 2.14 1.345 ;
        RECT 0.32 1.285 2.14 1.345 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.82 0.32 1.185 ;
        RECT 1.86 0.82 1.94 1.185 ;
        RECT 0.26 1.125 1.94 1.185 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 0.835 0.54 0.895 ;
        RECT 0.46 0.79 0.54 0.92 ;
        RECT 0.48 0.79 0.54 1.025 ;
        RECT 1.6 0.845 1.66 1.025 ;
        RECT 0.48 0.965 1.66 1.025 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.625 1.395 0.705 ;
        RECT 1.335 0.625 1.395 0.865 ;
        RECT 0.685 0.805 1.395 0.865 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.4 0.94 0.705 ;
        RECT 0.86 0.625 1.135 0.705 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END NAND4X2

MACRO DFFSRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX1 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.54 0.14 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.035 0.445 6.115 0.895 ;
        RECT 6.035 0.815 6.165 0.895 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.165 0.805 5.245 1.005 ;
        RECT 5.165 0.815 5.255 1.005 ;
        RECT 5.165 0.815 5.545 0.895 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.42 0.775 1.54 0.835 ;
        RECT 1.46 0.775 1.52 1.26 ;
        RECT 1.46 0.775 1.54 0.92 ;
        RECT 1.46 1.2 1.9 1.26 ;
        RECT 1.84 1.14 2.355 1.2 ;
        RECT 2.295 1.14 2.355 1.345 ;
        RECT 3.3 1.22 3.36 1.345 ;
        RECT 2.295 1.285 3.36 1.345 ;
        RECT 3.3 1.22 3.74 1.28 ;
        RECT 3.68 1.22 3.74 1.44 ;
        RECT 3.68 1.38 3.99 1.44 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 0.71 1.115 0.79 ;
        RECT 1.035 0.71 1.115 0.895 ;
        RECT 1.035 0.815 1.32 0.895 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END DFFSRHQX1

MACRO TLATNTSCAX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX3 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.415 0.9 3.475 1.29 ;
        RECT 3.46 0.52 3.52 0.96 ;
        RECT 3.46 0.6 3.54 0.73 ;
        RECT 3.415 0.9 3.885 0.96 ;
        RECT 3.825 0.9 3.885 1.29 ;
        RECT 3.87 0.52 3.93 0.66 ;
        RECT 3.46 0.6 3.93 0.66 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.765 0.925 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.6 0.515 0.925 ;
        RECT 0.46 0.45 0.54 0.73 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.035 0.525 0.175 0.895 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END TLATNTSCAX3

MACRO BUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX16 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.585 0.29 0.965 ;
        RECT 0.275 0.525 0.335 0.645 ;
        RECT 0.26 0.905 0.335 1.345 ;
        RECT 0.26 0.905 0.34 1.11 ;
        RECT 0.685 0.905 0.745 1.345 ;
        RECT 0.655 0.57 0.775 0.645 ;
        RECT 1.095 0.905 1.155 1.345 ;
        RECT 1.065 0.57 1.185 0.645 ;
        RECT 1.505 0.905 1.565 1.345 ;
        RECT 1.475 0.57 1.595 0.645 ;
        RECT 1.915 0.905 1.975 1.345 ;
        RECT 1.885 0.57 2.005 0.645 ;
        RECT 2.325 0.905 2.385 1.345 ;
        RECT 2.295 0.57 2.415 0.645 ;
        RECT 0.23 0.905 2.795 0.965 ;
        RECT 0.23 0.585 2.735 0.645 ;
        RECT 2.735 0.905 2.795 1.345 ;
        RECT 2.69 0.57 2.825 0.63 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.815 3.76 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END BUFX16

MACRO AOI33XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 0.29 0.865 0.41 ;
        RECT 1.04 1.11 1.1 1.265 ;
        RECT 0.805 0.35 1.51 0.41 ;
        RECT 1.45 0.35 1.51 1.3 ;
        RECT 1.04 1.11 1.51 1.17 ;
        RECT 1.45 1.17 1.54 1.3 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 1.1 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.51 1.14 0.99 ;
        RECT 1.06 0.51 1.16 0.63 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.51 1.34 1.01 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.54 0.35 ;
        RECT 0.48 0.27 0.56 0.7 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 1.1 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END AOI33XL

MACRO TLATSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRXL 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 1.005 0.73 ;
        RECT 0.925 0.49 1.005 1.22 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.02 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 0.98 3.54 1.185 ;
        RECT 3.59 0.815 3.67 1.06 ;
        RECT 3.46 0.98 3.67 1.06 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.2 0.815 2.63 0.895 ;
        RECT 2.435 0.815 2.63 0.965 ;
    END
  END RN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.61 1.94 1.11 ;
    END
  END G
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.815 1.6 1.06 ;
        RECT 1.265 0.96 1.6 1.06 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END TLATSRXL

MACRO MXI2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X8 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.06 0.405 2.12 1.425 ;
        RECT 2.06 0.98 2.14 1.11 ;
        RECT 2.47 0.98 2.53 1.425 ;
        RECT 2.44 0.435 2.56 0.495 ;
        RECT 2.85 0.435 2.97 0.51 ;
        RECT 2.88 0.98 2.94 1.425 ;
        RECT 2.91 0.435 2.97 1.04 ;
        RECT 2.06 0.98 3.35 1.04 ;
        RECT 3.29 0.39 3.35 0.51 ;
        RECT 2.515 0.45 3.35 0.51 ;
        RECT 3.29 0.98 3.35 1.425 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.705 1.34 1.205 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.645 0.54 1.025 ;
        RECT 0.46 0.645 0.66 0.92 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.34 1.11 ;
        RECT 0.28 0.99 0.36 1.205 ;
        RECT 0.76 0.865 0.84 1.205 ;
        RECT 0.28 1.125 0.84 1.205 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.6 0.06 ;
    END
  END VSS
END MXI2X8

MACRO CLKMX2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 0.365 1.525 0.485 ;
        RECT 1.465 1.045 1.525 1.435 ;
        RECT 1.5 0.425 1.56 1.105 ;
        RECT 1.5 0.6 1.74 0.66 ;
        RECT 1.66 0.6 1.74 0.73 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.22 0.815 1.3 1.215 ;
        RECT 1.22 0.815 1.4 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.635 0.54 1.035 ;
        RECT 0.44 0.955 0.62 1.035 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.34 1.215 ;
        RECT 0.72 0.93 0.8 1.215 ;
        RECT 0.26 1.135 0.8 1.215 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END CLKMX2X2

MACRO MX2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X6 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.61 0.295 1.67 0.415 ;
        RECT 1.635 0.83 1.695 1.395 ;
        RECT 1.655 0.355 1.715 0.88 ;
        RECT 1.655 0.6 1.74 0.88 ;
        RECT 2.02 0.235 2.08 0.66 ;
        RECT 2.045 0.6 2.105 1.395 ;
        RECT 1.655 0.6 2.47 0.66 ;
        RECT 2.41 0.485 2.47 0.985 ;
        RECT 2.43 0.235 2.49 0.545 ;
        RECT 2.455 0.925 2.515 1.395 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.675 1.34 1.175 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.615 0.66 0.995 ;
        RECT 0.46 0.79 0.66 0.995 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.915 0.36 1.11 ;
        RECT 0.76 0.915 0.84 1.175 ;
        RECT 0.28 1.095 0.84 1.175 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END MX2X6

MACRO MXI2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X6 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.03 0.29 2.09 0.76 ;
        RECT 2.03 0.86 2.09 1.48 ;
        RECT 2.03 0.7 2.32 0.76 ;
        RECT 2.26 0.7 2.32 0.92 ;
        RECT 2.26 0.79 2.34 0.92 ;
        RECT 2.03 0.86 2.34 0.92 ;
        RECT 2.44 0.29 2.5 1.48 ;
        RECT 2.26 0.79 2.91 0.85 ;
        RECT 2.805 0.63 2.865 0.85 ;
        RECT 2.85 0.29 2.91 0.69 ;
        RECT 2.85 0.79 2.91 1.48 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.76 1.34 1.26 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 1.1 ;
        RECT 0.59 0.73 0.67 0.92 ;
        RECT 0.46 0.79 0.67 0.92 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.34 1.11 ;
        RECT 0.3 1.05 0.36 1.26 ;
        RECT 0.77 0.96 0.83 1.26 ;
        RECT 0.3 1.2 0.83 1.26 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END MXI2X6

MACRO XOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.925 0.665 3.295 0.725 ;
        RECT 3.235 0.665 3.295 0.935 ;
        RECT 3.235 0.815 3.365 0.935 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.525 0.51 0.895 ;
        RECT 0.43 0.815 0.64 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.17 0.92 ;
        RECT 0.09 0.615 0.17 1.085 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.24 0.57 4.365 0.705 ;
        RECT 4.235 0.625 4.365 0.705 ;
        RECT 4.305 0.57 4.365 1.085 ;
        RECT 4.24 1.025 4.365 1.085 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
END XOR3X1

MACRO MDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.47 0.655 4.53 0.93 ;
        RECT 5.035 0.625 5.165 0.715 ;
        RECT 4.47 0.655 5.165 0.715 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.82 0.815 5.06 0.985 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.79 3.94 0.92 ;
        RECT 3.86 0.84 4.21 0.92 ;
        RECT 4.13 0.75 4.21 0.93 ;
    END
  END D0
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.69 0.34 1.19 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 1.075 ;
        RECT 0.525 0.54 0.585 0.85 ;
        RECT 1.005 0.54 1.065 1.075 ;
        RECT 0.46 1.015 1.065 1.075 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END MDFFHQX4

MACRO OAI211X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 1.17 0.685 1.45 ;
        RECT 1.07 0.38 1.13 0.5 ;
        RECT 1.06 1.17 1.14 1.45 ;
        RECT 1.11 0.44 1.17 1.23 ;
        RECT 0.625 1.17 1.17 1.23 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.9 0.14 1.11 ;
        RECT 0.21 0.76 0.29 1.085 ;
        RECT 0.06 0.9 0.29 1.085 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.64 0.54 0.72 ;
        RECT 0.46 0.64 0.54 1.07 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.79 0.74 1.07 ;
        RECT 0.71 0.64 0.79 0.895 ;
        RECT 0.64 0.79 0.79 0.895 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.41 0.97 0.54 ;
        RECT 0.89 0.41 0.97 0.84 ;
        RECT 0.89 0.76 1.01 0.84 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OAI211X1

MACRO TBUFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFXL 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.675 0.485 1.735 0.605 ;
        RECT 1.685 0.565 1.745 1.11 ;
        RECT 1.66 0.98 1.745 1.11 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.965 0.565 1.085 ;
        RECT 0.625 0.305 0.685 0.685 ;
        RECT 0.625 0.625 0.845 0.685 ;
        RECT 0.785 0.625 0.845 1.025 ;
        RECT 0.385 0.965 0.845 1.025 ;
        RECT 0.625 0.305 1.415 0.365 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.865 ;
        RECT 0.2 0.745 0.34 0.865 ;
        RECT 0.2 0.785 0.685 0.865 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END TBUFXL

MACRO DFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX1 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 0.73 ;
        RECT 0.88 0.495 0.94 1.455 ;
        RECT 0.92 0.435 0.98 0.555 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.29 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 0.755 1.965 0.96 ;
        RECT 1.795 0.805 2.17 0.96 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.04 0.815 1.365 1.06 ;
        RECT 1.04 0.935 1.375 1.06 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.435 0.625 4.655 0.815 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END DFFRX1

MACRO AND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.47 1.34 1.43 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.71 0.94 1.21 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.26 0.79 0.6 0.87 ;
        RECT 0.52 0.79 0.6 0.98 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.69 0.16 1.17 ;
        RECT 0.06 0.98 0.16 1.17 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END AND3X1

MACRO OAI222X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X2 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 1.155 0.685 1.275 ;
        RECT 1.685 1.155 1.745 1.275 ;
        RECT 2.415 0.415 2.475 0.555 ;
        RECT 2.52 1.155 2.58 1.275 ;
        RECT 2.825 0.415 2.885 0.555 ;
        RECT 2.415 0.495 3.32 0.555 ;
        RECT 3.26 0.495 3.32 1.215 ;
        RECT 0.625 1.155 3.32 1.215 ;
        RECT 3.26 0.6 3.34 0.73 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.845 0.335 1.055 ;
        RECT 0.86 0.79 0.94 1.055 ;
        RECT 0.275 0.995 0.94 1.055 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.42 0.835 1.54 0.895 ;
        RECT 1.46 0.79 1.54 1.055 ;
        RECT 2.08 0.845 2.14 1.055 ;
        RECT 1.46 0.995 2.14 1.055 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.845 2.32 1.055 ;
        RECT 2.86 0.79 2.92 1.055 ;
        RECT 2.26 0.995 2.92 1.055 ;
        RECT 2.86 0.79 2.94 0.92 ;
        RECT 2.86 0.79 2.98 0.85 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.675 0.65 0.895 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 0.655 2.76 0.895 ;
        RECT 2.42 0.775 2.76 0.895 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 0.655 1.98 0.735 ;
        RECT 1.835 0.655 1.98 0.895 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END OAI222X2

MACRO OAI33X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X4 0 0 ;
  SIZE 5.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.025 0.995 2.085 1.185 ;
        RECT 2.035 0.815 2.165 0.895 ;
        RECT 2.105 0.655 2.165 1.055 ;
        RECT 2.435 0.995 2.495 1.185 ;
        RECT 2.855 0.995 2.915 1.345 ;
        RECT 3.03 0.475 3.09 0.715 ;
        RECT 2.105 0.655 3.09 0.715 ;
        RECT 3.03 0.475 3.15 0.585 ;
        RECT 3.265 0.995 3.325 1.185 ;
        RECT 3.45 0.475 3.57 0.585 ;
        RECT 2.025 0.995 3.745 1.055 ;
        RECT 3.685 0.995 3.745 1.185 ;
        RECT 3.86 0.475 3.98 0.585 ;
        RECT 4.27 0.475 4.39 0.585 ;
        RECT 4.68 0.475 4.8 0.585 ;
        RECT 3.03 0.525 5.135 0.585 ;
        RECT 5.075 0.475 5.21 0.535 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.85 0.685 4.93 0.895 ;
        RECT 4.85 0.815 5.34 0.895 ;
    END
  END B0
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.14 0.815 3.64 0.895 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.25 0.815 1.74 0.895 ;
        RECT 1.66 0.655 1.74 0.92 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.265 0.815 2.765 0.895 ;
    END
  END A2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.655 0.94 0.92 ;
        RECT 0.495 0.84 0.94 0.92 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.01 0.685 4.165 0.895 ;
        RECT 4.01 0.815 4.455 0.895 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.8 0.06 ;
    END
  END VSS
END OAI33X4

MACRO MXI2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X4 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.75 0.835 1.81 1.35 ;
        RECT 1.905 0.43 1.965 0.895 ;
        RECT 1.795 0.815 1.965 0.895 ;
        RECT 1.75 0.835 2.22 0.895 ;
        RECT 2.16 0.835 2.22 1.35 ;
        RECT 1.77 0.43 2.36 0.49 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.45 0.64 1.53 1.13 ;
        RECT 1.45 0.8 1.54 1.13 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.64 0.71 0.92 ;
        RECT 0.63 0.64 0.71 0.97 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.965 0.34 1.11 ;
        RECT 0.81 0.925 0.87 1.13 ;
        RECT 0.28 1.07 0.87 1.13 ;
        RECT 1.13 0.595 1.19 1.045 ;
        RECT 0.81 0.985 1.19 1.045 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END MXI2X4

MACRO CLKAND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X4 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.135 0.425 1.195 0.565 ;
        RECT 1.235 0.945 1.295 1.335 ;
        RECT 1.545 0.425 1.605 0.565 ;
        RECT 1.235 0.945 1.74 1.005 ;
        RECT 1.135 0.505 1.72 0.565 ;
        RECT 1.66 0.505 1.72 1.335 ;
        RECT 1.66 0.79 1.74 1.335 ;
        RECT 1.645 0.945 1.74 1.335 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 0.815 0.765 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.625 0.565 0.715 ;
        RECT 0.285 0.635 0.875 0.715 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END CLKAND2X4

MACRO DFFSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX1 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.49 0.94 1.29 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.305 0.73 ;
        RECT 0.225 0.54 0.305 1.29 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.66 0.46 4.74 0.96 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.48 4.54 0.98 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.785 0.815 2.19 0.895 ;
        RECT 1.835 0.815 2.19 0.99 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END DFFSX1

MACRO FILL2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL2 0 0 ;
  SIZE 0.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.4 0.06 ;
    END
  END VSS
END FILL2

MACRO DFFNSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRXL 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.88 0.615 0.94 0.945 ;
        RECT 0.86 0.79 0.94 0.945 ;
        RECT 0.89 0.535 0.95 0.655 ;
        RECT 0.9 0.895 0.96 1.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.315 0.73 ;
        RECT 0.235 0.54 0.315 1.02 ;
    END
  END QN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.915 0.57 6.17 0.705 ;
        RECT 6.09 0.57 6.17 0.895 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.25 0.535 5.33 0.73 ;
        RECT 5.31 0.6 5.39 0.975 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 1.005 1.965 1.085 ;
        RECT 1.905 0.9 1.965 1.28 ;
        RECT 1.905 0.9 2.025 0.96 ;
        RECT 1.905 1.22 3.88 1.28 ;
        RECT 3.82 1.22 3.88 1.495 ;
        RECT 3.82 1.435 4.335 1.495 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.895 1.14 1.11 ;
        RECT 1.06 0.98 1.315 1.11 ;
        RECT 1.235 0.98 1.315 1.22 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.2 0.06 ;
    END
  END VSS
END DFFNSRXL

MACRO OAI211X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 1.005 0.76 1.345 ;
        RECT 1.36 1.005 1.42 1.345 ;
        RECT 1.94 0.655 2 1.065 ;
        RECT 1.99 1.005 2.05 1.345 ;
        RECT 0.7 1.005 2.165 1.065 ;
        RECT 2.4 1.025 2.46 1.345 ;
        RECT 2.795 0.525 2.855 0.715 ;
        RECT 1.94 0.655 2.855 0.715 ;
        RECT 2.81 1.025 2.87 1.345 ;
        RECT 3.015 0.445 3.075 0.585 ;
        RECT 1.99 1.025 3.28 1.085 ;
        RECT 3.22 1.025 3.28 1.345 ;
        RECT 3.425 0.445 3.485 0.585 ;
        RECT 2.795 0.525 3.485 0.585 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.605 0.815 1.375 0.895 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 0.66 0.34 0.72 ;
        RECT 0.26 0.66 0.34 0.92 ;
        RECT 0.305 0.655 1.685 0.715 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.93 0.79 3.355 0.87 ;
        RECT 3.06 0.79 3.14 0.92 ;
        RECT 3.275 0.76 3.355 0.88 ;
        RECT 3.06 0.79 3.355 0.88 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 0.815 2.6 0.895 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END OAI211X4

MACRO TLATNCAX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX8 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.24 0.54 3.3 1.395 ;
        RECT 3.24 0.6 3.34 1.01 ;
        RECT 3.65 0.95 3.71 1.395 ;
        RECT 3.62 0.57 3.74 0.63 ;
        RECT 4.06 0.95 4.12 1.395 ;
        RECT 4.03 0.57 4.15 0.645 ;
        RECT 3.695 0.585 4.53 0.645 ;
        RECT 3.24 0.95 4.53 1.01 ;
        RECT 4.47 0.525 4.53 1.395 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.81 0.66 1.15 ;
        RECT 0.58 1.005 0.775 1.15 ;
        RECT 0.535 1.07 0.775 1.15 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.355 0.75 0.435 1.085 ;
        RECT 0.19 1.005 0.435 1.085 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END TLATNCAX8

MACRO BUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX12 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.475 0.295 1.04 ;
        RECT 0.28 0.255 0.34 0.535 ;
        RECT 0.26 0.98 0.34 1.45 ;
        RECT 0.69 0.255 0.75 0.535 ;
        RECT 0.69 0.98 0.75 1.45 ;
        RECT 1.1 0.255 1.16 0.535 ;
        RECT 1.1 0.98 1.16 1.45 ;
        RECT 1.51 0.255 1.57 0.535 ;
        RECT 1.51 0.98 1.57 1.45 ;
        RECT 0.235 0.98 1.98 1.04 ;
        RECT 1.92 0.255 1.98 0.535 ;
        RECT 0.235 0.475 1.98 0.535 ;
        RECT 1.92 0.98 1.98 1.45 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.795 2.34 1.23 ;
        RECT 2.26 0.795 2.405 0.875 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END BUFX12

MACRO SEDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFX1 0 0 ;
  SIZE 7 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.635 0.54 3.695 0.705 ;
        RECT 3.635 0.625 3.82 0.705 ;
        RECT 3.76 0.625 3.82 1.095 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 0.49 1.94 0.61 ;
        RECT 1.86 0.49 1.94 0.99 ;
        RECT 1.86 0.91 1.98 0.99 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.66 0.79 6.88 0.98 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.62 3.34 1.12 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.98 2.34 1.12 ;
        RECT 2.365 0.725 2.445 1.06 ;
        RECT 2.26 0.98 2.445 1.06 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.54 0.815 0.88 0.935 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.38 0.655 0.44 0.895 ;
        RECT 0.235 0.815 0.44 0.895 ;
        RECT 0.885 0.335 0.945 0.715 ;
        RECT 0.38 0.655 1.04 0.715 ;
        RECT 0.98 0.655 1.04 0.78 ;
        RECT 0.885 0.335 1.52 0.395 ;
        RECT 1.46 0.335 1.52 0.91 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7 0.06 ;
    END
  END VSS
END SEDFFX1

MACRO OAI33X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X2 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.03 1.005 3.165 1.085 ;
        RECT 3.97 0.945 4.03 1.065 ;
        RECT 2.84 1.005 4.03 1.065 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 0.995 2.235 1.055 ;
        RECT 2.035 0.995 2.235 1.085 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 0.845 2.74 1.11 ;
        RECT 2.66 0.98 2.74 1.11 ;
        RECT 2.68 0.845 3.87 0.905 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.485 0.815 1.935 0.875 ;
        RECT 1.635 0.815 1.935 0.895 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.46 0.685 2.54 0.92 ;
        RECT 2.46 0.685 3.71 0.745 ;
    END
  END B2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.625 0.565 0.705 ;
        RECT 0.325 0.645 1.5 0.705 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.475 0.415 2.595 0.515 ;
        RECT 2.435 0.435 2.595 0.515 ;
        RECT 2.535 0.415 2.595 0.585 ;
        RECT 2.915 0.415 3.035 0.585 ;
        RECT 3.355 0.415 3.475 0.585 ;
        RECT 3.795 0.415 3.87 0.585 ;
        RECT 2.535 0.525 3.87 0.585 ;
        RECT 3.795 0.415 3.915 0.475 ;
        RECT 4.13 0.575 4.19 1.27 ;
        RECT 0.835 1.21 4.19 1.27 ;
        RECT 4.19 0.445 4.25 0.635 ;
        RECT 3.81 0.575 4.25 0.635 ;
        RECT 4.235 0.385 4.295 0.505 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END OAI33X2

MACRO EDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX2 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.79 3.125 0.92 ;
        RECT 3.045 0.55 3.125 1.14 ;
        RECT 3.045 0.55 3.165 0.63 ;
        RECT 3.045 1.06 3.175 1.14 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.79 0.28 3.85 0.98 ;
        RECT 4.11 0.6 4.17 0.8 ;
        RECT 3.79 0.28 4.295 0.34 ;
        RECT 4.235 0.28 4.295 0.66 ;
        RECT 4.11 0.6 4.94 0.66 ;
        RECT 4.86 0.6 4.94 0.73 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.76 4.54 1.03 ;
        RECT 4.45 0.76 4.76 0.84 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.745 0.31 1.085 ;
        RECT 0.235 1.005 0.425 1.13 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.2 0.06 ;
    END
  END VSS
END EDFFHQX2

MACRO AND4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 1.005 1.565 1.085 ;
        RECT 1.425 0.505 1.485 0.625 ;
        RECT 1.425 0.565 1.565 0.625 ;
        RECT 1.505 0.565 1.565 1.47 ;
        RECT 1.47 1.005 1.565 1.47 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.775 1.165 0.92 ;
        RECT 1.085 0.775 1.165 1.25 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.725 0.74 1.225 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.98 0.54 1.205 ;
        RECT 0.48 0.725 0.56 1.06 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 0.76 0.34 0.84 ;
        RECT 0.26 0.725 0.34 1.185 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END AND4X1

MACRO CLKMX2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X8 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2 0.53 2.12 0.59 ;
        RECT 2.035 0.99 2.095 1.435 ;
        RECT 2.06 0.53 2.12 1.11 ;
        RECT 2.06 0.98 2.14 1.11 ;
        RECT 2.445 0.99 2.505 1.435 ;
        RECT 2.415 0.54 2.535 0.6 ;
        RECT 2.855 0.99 2.915 1.435 ;
        RECT 2.825 0.54 2.945 0.615 ;
        RECT 2.49 0.555 3.325 0.615 ;
        RECT 2.035 0.99 3.325 1.05 ;
        RECT 3.265 0.495 3.325 1.435 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 0.85 1.74 0.93 ;
        RECT 1.66 0.85 1.74 1.19 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.715 0.8 1.085 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.955 0.535 1.11 ;
        RECT 0.475 0.955 0.535 1.245 ;
        RECT 0.9 0.865 0.96 1.245 ;
        RECT 0.475 1.185 0.96 1.245 ;
        RECT 0.9 0.865 1.02 0.925 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END CLKMX2X8

MACRO XNOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.2 0.54 ;
        RECT 0.14 0.41 0.2 1.335 ;
        RECT 0.235 0.35 0.295 0.47 ;
        RECT 0.06 0.41 0.295 0.47 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.19 0.815 1.57 0.895 ;
        RECT 1.49 0.735 1.61 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 0.97 ;
        RECT 0.53 0.54 0.61 0.87 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END XNOR2X1

MACRO AOI22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X4 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.695 0.445 0.815 0.505 ;
        RECT 1.315 0.445 1.435 0.525 ;
        RECT 1.74 0.465 1.8 0.895 ;
        RECT 1.74 0.815 1.965 0.895 ;
        RECT 1.96 0.835 2.02 1.115 ;
        RECT 2.135 0.445 2.255 0.525 ;
        RECT 2.37 0.995 2.43 1.115 ;
        RECT 0.765 0.465 2.715 0.525 ;
        RECT 2.78 0.995 2.84 1.115 ;
        RECT 2.665 0.445 2.875 0.505 ;
        RECT 1.96 0.995 3.25 1.055 ;
        RECT 3.19 0.995 3.25 1.115 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.21 0.815 2.945 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 0.815 1.36 0.895 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.215 0.655 1.64 0.715 ;
        RECT 1.46 0.655 1.54 0.92 ;
        RECT 1.58 0.625 1.64 0.745 ;
        RECT 1.46 0.655 1.64 0.745 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 0.625 2.165 0.705 ;
        RECT 1.9 0.645 3.355 0.705 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.6 0.06 ;
    END
  END VSS
END AOI22X4

MACRO SMDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX4 0 0 ;
  SIZE 6.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 0.645 5.66 0.99 ;
        RECT 5.6 0.645 6.39 0.705 ;
        RECT 6.235 0.625 6.365 0.705 ;
        RECT 6.33 0.645 6.39 0.765 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.93 0.805 6.165 1.085 ;
        RECT 5.93 0.805 6.23 0.885 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.455 5.34 0.955 ;
    END
  END D0
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.455 5.14 0.955 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.025 0.585 4.105 0.92 ;
        RECT 3.86 0.79 4.105 0.92 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.42 0.34 0.92 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.53 0.535 0.59 1.05 ;
        RECT 0.46 0.79 0.59 1.05 ;
        RECT 0.895 0.65 0.955 1.05 ;
        RECT 0.94 0.535 1 0.71 ;
        RECT 0.46 0.99 1.13 1.05 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.8 0.06 ;
    END
  END VSS
END SMDFFHQX4

MACRO BUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX3 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 0.48 0.235 0.62 ;
        RECT 0.215 1.05 0.275 1.44 ;
        RECT 0.26 0.56 0.32 1.11 ;
        RECT 0.26 0.98 0.34 1.11 ;
        RECT 0.54 0.405 0.6 0.62 ;
        RECT 0.175 0.56 0.6 0.62 ;
        RECT 0.215 1.05 0.685 1.11 ;
        RECT 0.585 0.345 0.645 0.465 ;
        RECT 0.625 1.05 0.685 1.44 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.72 0.94 1.22 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END BUFX3

MACRO TLATNCAX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX20 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.355 4.52 0.92 ;
        RECT 4.49 0.785 4.55 1.405 ;
        RECT 4.87 0.355 4.93 0.845 ;
        RECT 4.9 0.785 4.96 1.405 ;
        RECT 5.235 0.6 5.295 0.845 ;
        RECT 5.28 0.355 5.34 0.66 ;
        RECT 5.31 0.785 5.37 1.405 ;
        RECT 5.69 0.355 5.75 0.845 ;
        RECT 5.72 0.785 5.78 1.405 ;
        RECT 6.055 0.625 6.115 0.845 ;
        RECT 6.1 0.355 6.16 0.685 ;
        RECT 6.13 0.785 6.19 1.405 ;
        RECT 6.51 0.355 6.57 0.845 ;
        RECT 6.54 0.785 6.6 1.405 ;
        RECT 6.875 0.6 6.935 0.845 ;
        RECT 6.92 0.355 6.98 0.66 ;
        RECT 6.95 0.785 7.01 1.405 ;
        RECT 7.33 0.355 7.39 0.845 ;
        RECT 7.36 0.785 7.42 1.405 ;
        RECT 7.695 0.6 7.755 0.845 ;
        RECT 4.46 0.785 7.83 0.845 ;
        RECT 7.74 0.355 7.8 0.66 ;
        RECT 7.77 0.785 7.83 1.4 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8 0.06 ;
    END
  END VSS
END TLATNCAX20

MACRO AOI22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X2 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.165 0.415 1.225 0.895 ;
        RECT 1.035 0.815 1.225 0.895 ;
        RECT 1.035 0.835 1.49 0.895 ;
        RECT 1.43 0.835 1.49 1.165 ;
        RECT 0.71 0.415 1.685 0.475 ;
        RECT 1.84 0.995 1.9 1.165 ;
        RECT 1.43 1.105 1.9 1.165 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 0.715 0.745 0.96 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.74 1.74 1.03 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 0.58 1.56 0.715 ;
        RECT 1.325 0.655 1.56 0.715 ;
        RECT 1.5 0.58 1.96 0.64 ;
        RECT 1.84 0.58 1.96 0.895 ;
        RECT 1.84 0.815 2.165 0.895 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.56 0.705 ;
        RECT 0.48 0.575 0.92 0.655 ;
        RECT 0.84 0.635 1.065 0.715 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END AOI22X2

MACRO MXI3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3X4 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.015 0.965 2.075 1.35 ;
        RECT 2.06 0.79 2.12 1.025 ;
        RECT 2.06 0.79 2.14 0.92 ;
        RECT 2.06 0.86 2.485 0.92 ;
        RECT 2.425 0.47 2.485 1.35 ;
        RECT 2.02 0.47 2.61 0.53 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 0.645 3.06 1.015 ;
        RECT 3.235 0.625 3.325 0.765 ;
        RECT 3.235 0.625 3.365 0.705 ;
        RECT 3 0.645 3.71 0.705 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.635 0.805 3.77 0.945 ;
        RECT 3.33 0.865 3.77 0.945 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.63 2.74 1.13 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.79 0.825 0.85 ;
        RECT 0.765 0.77 1.09 0.83 ;
        RECT 1.06 0.6 1.14 0.77 ;
        RECT 1.03 0.685 1.14 0.77 ;
        RECT 1.03 0.71 1.41 0.77 ;
        RECT 1.35 0.71 1.41 0.955 ;
        RECT 1.35 0.895 1.47 0.955 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.06 0.46 0.255 0.54 ;
        RECT 0.175 0.46 0.255 0.795 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END MXI3X4

MACRO TLATNCAX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.52 0.74 0.73 ;
        RECT 0.67 0.68 0.75 1.02 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.615 0.67 2.695 1.055 ;
        RECT 2.615 0.815 2.81 0.935 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.38 0.65 0.46 1.02 ;
        RECT 0.46 0.6 0.54 0.73 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END TLATNCAX2

MACRO OAI2BB1X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.61 0.23 1.17 ;
        RECT 0.06 0.98 0.23 1.17 ;
        RECT 0.39 1.11 0.45 1.48 ;
        RECT 0.595 0.53 0.655 0.67 ;
        RECT 0.17 0.61 0.655 0.67 ;
        RECT 0.06 1.11 0.86 1.17 ;
        RECT 0.8 1.11 0.86 1.48 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.77 0.54 0.92 ;
        RECT 0.33 0.77 0.92 0.85 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.02 0.625 1.165 0.705 ;
        RECT 1.085 0.625 1.165 0.85 ;
        RECT 1.085 0.77 1.375 0.85 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.825 1.715 1.25 ;
        RECT 1.66 1.17 1.74 1.3 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OAI2BB1X2

MACRO MXI2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X2 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.845 0.46 1.905 0.6 ;
        RECT 1.86 0.54 1.92 1.335 ;
        RECT 1.86 0.6 1.94 0.73 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.7 1.54 1.115 ;
        RECT 1.46 0.7 1.625 0.92 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.7 0.765 0.955 ;
        RECT 0.44 0.79 0.765 0.955 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.95 0.34 1.11 ;
        RECT 0.865 0.84 0.925 1.115 ;
        RECT 0.28 1.055 0.925 1.115 ;
        RECT 1.14 0.7 1.2 0.9 ;
        RECT 0.865 0.84 1.2 0.9 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END MXI2X2

MACRO FILL64
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL64 0 0 ;
  SIZE 12.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 12.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 12.8 0.06 ;
    END
  END VSS
END FILL64

MACRO SMDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX1 0 0 ;
  SIZE 6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.145 0.73 ;
        RECT 0.085 0.54 0.145 1.34 ;
    END
  END Q
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5 0.77 5.06 1.04 ;
        RECT 5.075 0.645 5.135 0.83 ;
        RECT 5 0.77 5.135 0.83 ;
        RECT 5.235 0.625 5.365 0.705 ;
        RECT 5.075 0.645 5.79 0.705 ;
        RECT 5.73 0.645 5.79 0.765 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.33 0.805 5.63 0.925 ;
        RECT 5.55 0.805 5.63 1.085 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.66 0.485 4.74 0.985 ;
    END
  END D0
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.6 4.54 1.1 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 0.585 3.54 0.82 ;
        RECT 3.535 0.6 3.615 1.01 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.92 0.34 1.11 ;
        RECT 0.43 0.78 0.51 1 ;
        RECT 0.26 0.92 0.51 1 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6 0.06 ;
    END
  END VSS
END SMDFFHQX1

MACRO TLATSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.275 0.5 4.335 0.62 ;
        RECT 4.275 0.875 4.335 1.345 ;
        RECT 4.32 0.56 4.38 0.935 ;
        RECT 4.32 0.79 4.54 0.92 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.455 0.415 3.515 0.535 ;
        RECT 3.455 0.85 3.515 1.345 ;
        RECT 3.475 0.475 3.535 0.91 ;
        RECT 3.475 0.625 3.765 0.685 ;
        RECT 3.635 0.625 3.765 0.705 ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 0.795 3.115 1.125 ;
        RECT 3.035 0.795 3.155 1.085 ;
        RECT 3.035 1.005 3.285 1.085 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.565 0.905 1.94 0.985 ;
        RECT 1.86 0.905 1.94 1.11 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.66 0.7 0.92 ;
        RECT 0.62 0.66 0.7 1 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.53 2.34 1.03 ;
    END
  END G
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END TLATSRX2

MACRO INVX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX20 0 0 ;
  SIZE 3.80 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.535 0.72 3.615 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.72 0.15 0.87 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.80 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.80 0.06 ;
    END
  END VSS
END INVX20

MACRO AOI32X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.64 0.335 2.7 0.895 ;
        RECT 2.64 0.815 2.965 0.895 ;
        RECT 2.87 0.815 2.965 1.115 ;
        RECT 3.28 0.995 3.34 1.115 ;
        RECT 3.69 0.995 3.75 1.115 ;
        RECT 0.835 0.335 3.845 0.395 ;
        RECT 2.87 0.995 4.16 1.055 ;
        RECT 4.1 0.995 4.16 1.115 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.855 0.815 1.165 0.895 ;
        RECT 1.11 0.835 1.17 0.985 ;
        RECT 1.855 0.815 1.915 0.985 ;
        RECT 1.11 0.925 1.915 0.985 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.12 0.815 3.855 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.655 0.74 0.92 ;
        RECT 0.535 0.655 1.33 0.715 ;
        RECT 1.27 0.655 1.33 0.825 ;
        RECT 1.675 0.655 1.735 0.825 ;
        RECT 1.27 0.765 1.735 0.825 ;
        RECT 1.675 0.655 2.32 0.715 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.375 0.495 0.435 0.695 ;
        RECT 1.43 0.495 1.55 0.665 ;
        RECT 0.375 0.495 2.52 0.555 ;
        RECT 2.42 0.655 2.54 0.715 ;
        RECT 2.46 0.495 2.52 0.73 ;
        RECT 2.46 0.6 2.54 0.73 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.8 0.625 3.165 0.705 ;
        RECT 2.8 0.645 4.265 0.705 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END AOI32X4

MACRO SDFFQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.54 0.14 1.34 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.49 0.745 3.55 1.005 ;
        RECT 3.515 0.645 3.575 0.805 ;
        RECT 3.685 0.585 3.745 0.705 ;
        RECT 3.685 0.625 4.165 0.705 ;
        RECT 3.515 0.645 4.165 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.835 0.805 3.965 1.01 ;
        RECT 3.835 0.805 4.21 0.885 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 0.625 3.23 0.705 ;
        RECT 3.15 0.62 3.23 1.005 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.92 0.34 1.115 ;
        RECT 0.425 0.78 0.505 1 ;
        RECT 0.26 0.92 0.505 1 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END SDFFQX1

MACRO INVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX4 0 0 ;
  SIZE 1.00 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.87 0.63 0.95 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.72 0.15 0.87 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.00 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.00 0.06 ;
    END
  END VSS
END INVX4

MACRO CLKMX2X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X12 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.54 0.415 1.6 0.535 ;
        RECT 1.54 0.475 1.695 0.535 ;
        RECT 1.635 0.475 1.695 1.48 ;
        RECT 1.635 0.79 1.74 0.92 ;
        RECT 2 0.3 2.06 0.85 ;
        RECT 2.045 0.79 2.105 1.48 ;
        RECT 2.41 0.3 2.47 0.85 ;
        RECT 2.455 0.79 2.515 1.48 ;
        RECT 2.82 0.3 2.88 0.85 ;
        RECT 2.865 0.79 2.925 1.48 ;
        RECT 1.635 0.79 3.29 0.85 ;
        RECT 3.23 0.3 3.29 0.98 ;
        RECT 3.275 0.92 3.335 1.48 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.225 0.99 1.305 1.26 ;
        RECT 1.26 0.795 1.34 1.11 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.68 0.56 1.08 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.92 0.34 1.26 ;
        RECT 0.66 1.035 0.74 1.26 ;
        RECT 0.26 1.18 0.74 1.26 ;
        RECT 0.66 1.035 0.805 1.115 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END CLKMX2X12

MACRO DFFSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRXL 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.945 0.73 ;
        RECT 0.885 0.575 0.945 1.315 ;
        RECT 0.94 0.515 1 0.635 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.315 0.73 ;
        RECT 0.235 0.54 0.315 1.02 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.755 6.34 1.255 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.66 0.485 5.74 0.925 ;
        RECT 5.66 0.79 5.8 0.925 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 0.625 3.165 0.765 ;
        RECT 3.105 0.3 3.165 0.765 ;
        RECT 2.04 0.705 3.165 0.765 ;
        RECT 3.105 0.3 3.805 0.36 ;
        RECT 3.745 0.3 3.805 0.86 ;
        RECT 3.745 0.8 4.605 0.86 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.195 0.9 1.365 1.16 ;
        RECT 1.045 1.005 1.365 1.16 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END DFFSRXL

MACRO EDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX8 0 0 ;
  SIZE 6.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.03 0.54 3.09 0.66 ;
        RECT 3.08 0.6 3.14 1.025 ;
        RECT 3.06 0.79 3.14 1.025 ;
        RECT 3.5 0.54 3.56 0.66 ;
        RECT 3.97 0.54 4.03 0.66 ;
        RECT 2.995 0.965 4.345 1.025 ;
        RECT 4.44 0.54 4.5 0.66 ;
        RECT 3.03 0.6 4.5 0.66 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.595 0.325 5.655 0.895 ;
        RECT 5.595 0.325 6.1 0.385 ;
        RECT 6.04 0.325 6.1 0.705 ;
        RECT 5.915 0.645 6.565 0.705 ;
        RECT 6.245 0.625 6.565 0.715 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.075 0.815 6.575 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.76 0.34 1.26 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.8 0.06 ;
    END
  END VSS
END EDFFHQX8

MACRO MXI3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3X2 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.06 0.57 2.14 1.335 ;
        RECT 2.05 0.57 2.17 0.65 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.635 0.84 2.695 0.96 ;
        RECT 2.69 0.49 2.75 0.9 ;
        RECT 2.9 0.49 2.96 0.68 ;
        RECT 2.69 0.49 3.555 0.55 ;
        RECT 3.435 0.49 3.555 0.705 ;
        RECT 3.435 0.625 3.565 0.705 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.255 0.65 3.335 0.955 ;
        RECT 3.06 0.79 3.335 0.955 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.79 2.34 0.92 ;
        RECT 2.295 0.455 2.375 0.87 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.72 0.88 0.78 1.065 ;
        RECT 0.835 1.005 0.965 1.085 ;
        RECT 1.22 0.71 1.28 1.065 ;
        RECT 1.485 0.87 1.545 1.065 ;
        RECT 0.72 1.005 1.545 1.065 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.98 0.14 1.11 ;
        RECT 0.18 0.73 0.26 1.06 ;
        RECT 0.06 0.98 0.26 1.06 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END MXI3X2

MACRO MX2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.48 0.37 1.54 1.415 ;
        RECT 1.48 0.98 1.74 1.11 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.72 1.365 1.09 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.61 0.635 1.015 ;
        RECT 0.46 0.79 0.635 1.015 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.34 1.195 ;
        RECT 0.735 0.835 0.815 1.195 ;
        RECT 0.26 1.115 0.815 1.195 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END MX2X1

MACRO SEDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX4 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.07 0.645 7.13 0.89 ;
        RECT 7.01 0.83 7.13 0.89 ;
        RECT 7.635 0.625 7.97 0.705 ;
        RECT 7.07 0.645 7.97 0.705 ;
        RECT 7.91 0.625 7.97 0.745 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.39 0.805 7.565 0.965 ;
        RECT 7.39 0.805 7.81 0.885 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.415 0.695 6.495 0.94 ;
        RECT 6.415 0.815 6.75 0.94 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.71 5.34 1.21 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.835 0.775 5.16 0.895 ;
        RECT 5.08 0.71 5.16 0.965 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.54 0.335 1.35 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.26 0.67 0.745 0.73 ;
        RECT 0.685 0.54 0.745 1.35 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.2 0.06 ;
    END
  END VSS
END SEDFFHQX4

MACRO MXI4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.835 0.775 2.895 1.315 ;
        RECT 4.625 1.095 4.685 1.315 ;
        RECT 2.835 1.255 4.685 1.315 ;
        RECT 4.835 0.815 4.965 0.895 ;
        RECT 4.905 0.815 4.965 1.155 ;
        RECT 4.625 1.095 4.965 1.155 ;
        RECT 4.835 0.815 5.205 0.875 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.08 0.375 4.14 0.645 ;
        RECT 4.14 0.585 4.2 0.995 ;
        RECT 4.08 0.935 4.2 0.995 ;
        RECT 4.46 0.585 4.54 0.73 ;
        RECT 4.48 0.585 4.54 0.995 ;
        RECT 4.48 0.935 4.67 0.995 ;
        RECT 4.78 0.375 4.84 0.645 ;
        RECT 4.08 0.585 4.84 0.645 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.445 0.75 2.525 1.1 ;
        RECT 2.46 0.98 2.575 1.2 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.68 0.72 1.76 1.2 ;
        RECT 1.66 0.98 1.76 1.2 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.98 1.54 1.2 ;
        RECT 1.48 0.72 1.56 1.1 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.865 0.58 1.205 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.685 0.34 0.92 ;
        RECT 0.26 0.685 0.89 0.765 ;
        RECT 0.81 0.685 0.89 0.94 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END MXI4X4

MACRO DLY1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY1X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.52 1.495 0.66 ;
        RECT 1.435 0.9 1.495 1.29 ;
        RECT 1.46 0.6 1.52 0.96 ;
        RECT 1.46 0.79 1.54 0.96 ;
        RECT 1.435 0.9 1.905 0.96 ;
        RECT 1.845 0.52 1.905 0.66 ;
        RECT 1.435 0.6 1.905 0.66 ;
        RECT 1.845 0.9 1.905 1.29 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.775 0.315 1.145 ;
        RECT 0.235 0.775 0.445 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END DLY1X4

MACRO SDFFSRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX2 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.54 0.42 0.8 ;
        RECT 0.4 0.74 0.46 1.09 ;
        RECT 0.445 1.03 0.505 1.3 ;
        RECT 0.445 1.17 0.54 1.3 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7 0.655 7.06 0.935 ;
        RECT 7 0.655 7.92 0.715 ;
        RECT 7.86 0.715 7.94 0.92 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.38 0.85 7.76 0.93 ;
        RECT 7.435 0.815 7.76 1.015 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.66 0.5 6.74 1 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.48 0.66 6.56 0.895 ;
        RECT 6.215 0.815 6.56 0.895 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.815 1.78 0.895 ;
        RECT 1.72 0.815 1.78 1 ;
        RECT 1.72 0.94 2.76 1 ;
        RECT 2.7 0.94 2.76 1.35 ;
        RECT 3.5 1.155 3.56 1.35 ;
        RECT 2.7 1.29 3.56 1.35 ;
        RECT 3.5 1.155 3.94 1.215 ;
        RECT 3.88 1.155 3.94 1.34 ;
        RECT 3.88 1.28 4.64 1.34 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.75 1.34 1 ;
        RECT 1.205 0.75 1.535 0.83 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.2 0.06 ;
    END
  END VSS
END SDFFSRHQX2

MACRO XOR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.2 0.73 ;
        RECT 0.12 0.44 0.2 1.18 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.875 0.815 0.935 0.935 ;
        RECT 1.035 0.815 1.165 0.895 ;
        RECT 1.13 0.8 1.25 0.875 ;
        RECT 0.875 0.815 1.54 0.875 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.98 0.54 1.25 ;
        RECT 0.535 0.825 0.615 1.06 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END XOR2XL

MACRO SEDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX1 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.6 3.34 0.73 ;
        RECT 3.485 0.67 3.545 1.29 ;
        RECT 3.545 0.54 3.605 0.73 ;
        RECT 3.26 0.67 3.605 0.73 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.61 6.34 1.11 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.705 0.68 2.825 0.895 ;
        RECT 2.705 0.815 2.975 0.895 ;
        RECT 2.835 0.815 2.975 0.99 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.54 0.625 1.805 0.705 ;
        RECT 1.725 0.625 1.805 0.94 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.475 0.655 0.555 0.97 ;
        RECT 0.475 0.79 0.74 0.97 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.365 0.705 ;
        RECT 0.315 0.495 0.375 0.685 ;
        RECT 0.315 0.495 0.96 0.555 ;
        RECT 0.9 0.495 0.96 0.695 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END SEDFFHQX1

MACRO TLATNXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNXL 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.405 3.14 1.02 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.405 2.34 1.385 ;
        RECT 2.26 1.265 2.355 1.385 ;
    END
  END QN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.06 0.76 2.14 1.26 ;
    END
  END GN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.955 0.34 1.12 ;
        RECT 0.4 0.76 0.48 1.11 ;
        RECT 0.26 0.955 0.48 1.11 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END TLATNXL

MACRO OAI2BB2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2XL 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 1.15 1.765 1.275 ;
        RECT 1.555 1.215 1.765 1.275 ;
        RECT 1.84 0.355 1.9 1.21 ;
        RECT 1.635 1.15 1.9 1.21 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2 0.65 2.08 1.04 ;
        RECT 2.06 0.6 2.14 0.73 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.55 1.74 1.05 ;
    END
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.59 0.54 1.09 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.5 0.34 1 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END OAI2BB2XL

MACRO OR4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.37 1.54 1.315 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 0.73 ;
        RECT 0.675 0.65 0.755 1.085 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.63 0.56 1.11 ;
        RECT 0.46 0.98 0.56 1.11 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.59 1.2 0.73 ;
        RECT 1.12 0.59 1.2 1.03 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END OR4XL

MACRO FILL8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL8 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END FILL8

MACRO DFFQXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQXL 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.495 0.14 1.31 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.755 0.845 2.965 1.185 ;
        RECT 2.73 1.105 2.965 1.185 ;
        RECT 2.755 0.845 2.97 0.925 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.85 0.485 1.185 ;
        RECT 0.24 0.98 0.485 1.185 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END DFFQXL

MACRO AND2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 0.73 ;
        RECT 0.87 0.53 0.94 1.235 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 0.945 0.705 1.25 ;
        RECT 0.66 1.17 0.74 1.41 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 1.025 ;
        RECT 0.285 0.75 0.365 0.87 ;
        RECT 0.06 0.79 0.365 0.87 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END AND2XL

MACRO CLKBUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX3 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 0.48 0.235 0.62 ;
        RECT 0.215 1.05 0.275 1.44 ;
        RECT 0.26 0.56 0.32 1.11 ;
        RECT 0.26 0.98 0.34 1.11 ;
        RECT 0.54 0.405 0.6 0.62 ;
        RECT 0.175 0.56 0.6 0.62 ;
        RECT 0.215 1.05 0.685 1.11 ;
        RECT 0.585 0.345 0.645 0.465 ;
        RECT 0.625 1.05 0.685 1.44 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.72 0.94 1.22 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END CLKBUFX3

MACRO DFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRXL 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.57 0.94 0.98 ;
        RECT 0.88 0.9 0.96 1.17 ;
        RECT 0.895 0.525 0.975 0.645 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.02 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.41 4.34 0.54 ;
        RECT 4.29 0.46 4.37 0.88 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.38 4.14 0.83 ;
        RECT 4.06 0.75 4.19 0.83 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.93 1.14 1.3 ;
        RECT 1.22 0.89 1.3 1.01 ;
        RECT 1.06 0.93 1.3 1.01 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END DFFTRXL

MACRO OR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X2 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.765 0.385 0.825 0.505 ;
        RECT 0.765 0.905 0.825 1.375 ;
        RECT 0.765 0.445 0.92 0.505 ;
        RECT 0.86 0.445 0.92 0.965 ;
        RECT 0.765 0.905 0.92 0.965 ;
        RECT 0.86 0.6 0.94 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 0.765 0.49 1.155 ;
        RECT 0.41 0.815 0.515 1.155 ;
        RECT 0.41 0.815 0.6 0.895 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.07 0.46 0.15 0.9 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OR2X2

MACRO DLY2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY2X4 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.06 0.6 2.14 1.075 ;
        RECT 2.035 0.84 2.14 1.075 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.365 0.495 0.425 1.335 ;
        RECT 0.365 0.6 0.54 0.73 ;
        RECT 0.365 0.6 0.79 0.66 ;
        RECT 0.73 0.415 0.79 1.175 ;
        RECT 0.775 0.355 0.835 0.475 ;
        RECT 0.775 1.115 0.835 1.335 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END DLY2X4

MACRO NAND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1 0 0 ;
  SIZE 0.60 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.475 0.76 0.555 0.9 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.095 0.805 0.215 0.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 0.615 0.375 0.745 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.60 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.60 0.06 ;
    END
  END VSS
END NAND2X1

MACRO MXI4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X2 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.605 0.565 4.725 0.645 ;
        RECT 4.645 0.565 4.725 1.025 ;
        RECT 4.645 0.79 4.74 0.92 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 1.005 1.92 1.25 ;
    END
  END C
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.65 0.345 0.92 ;
        RECT 0.26 0.65 0.73 0.73 ;
        RECT 0.65 0.65 0.73 0.86 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.15 1.005 1.365 1.25 ;
        RECT 1.15 1.015 1.485 1.25 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.83 0.54 1.14 ;
        RECT 0.46 0.96 0.73 1.04 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.305 0.875 3.365 1.315 ;
        RECT 3.39 0.79 3.45 0.935 ;
        RECT 3.305 0.875 3.45 0.935 ;
        RECT 4.96 0.835 5.02 1.315 ;
        RECT 3.305 1.255 5.02 1.315 ;
        RECT 5.035 0.765 5.165 0.895 ;
        RECT 4.96 0.835 5.165 0.895 ;
    END
  END S1
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.62 2.94 1.12 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END MXI4X2

MACRO AOI32X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X2 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.505 0.435 1.565 1.085 ;
        RECT 1.435 1.005 1.565 1.085 ;
        RECT 1.435 1.005 1.79 1.065 ;
        RECT 1.73 1.005 1.79 1.225 ;
        RECT 0.815 0.435 2.025 0.495 ;
        RECT 1.73 1.105 2.2 1.165 ;
        RECT 2.14 1.105 2.2 1.225 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.52 0.915 0.6 1.085 ;
        RECT 0.435 1.005 0.6 1.085 ;
        RECT 0.52 0.915 0.855 0.995 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.52 0.755 1.14 0.815 ;
        RECT 1.06 0.755 1.14 0.92 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.89 0.875 2.34 1.005 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.595 0.42 0.82 ;
        RECT 0.36 0.595 1.34 0.655 ;
        RECT 1.26 0.595 1.34 0.82 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.665 0.625 1.79 0.8 ;
        RECT 1.665 0.625 2.535 0.705 ;
        RECT 2.415 0.625 2.535 0.8 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END AOI32X2

MACRO DFFNSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX2 0 0 ;
  SIZE 7 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.355 0.54 6.435 1.06 ;
        RECT 6.355 0.98 6.54 1.06 ;
        RECT 6.46 0.98 6.54 1.11 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.86 0.54 5.94 1.11 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.78 0.54 1.26 ;
        RECT 0.46 0.98 0.56 1.26 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 0.575 3.025 0.92 ;
        RECT 2.945 0.73 3.14 0.92 ;
        RECT 3.06 0.73 3.14 0.96 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.585 0.575 2.665 0.895 ;
        RECT 2.585 0.815 2.845 0.895 ;
    END
  END SN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.78 0.34 0.92 ;
        RECT 0.28 0.79 0.36 1.26 ;
    END
  END CKN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7 0.06 ;
    END
  END VSS
END DFFNSRX2

MACRO OR3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X4 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.905 0.91 0.965 1.46 ;
        RECT 0.915 0.4 1.035 0.46 ;
        RECT 0.985 0.42 1.49 0.48 ;
        RECT 1.315 1.07 1.375 1.46 ;
        RECT 0.905 0.91 1.49 0.97 ;
        RECT 1.37 0.36 1.43 0.48 ;
        RECT 1.43 0.42 1.49 1.13 ;
        RECT 1.315 1.07 1.49 1.13 ;
        RECT 1.43 0.6 1.74 0.66 ;
        RECT 1.66 0.6 1.74 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.74 0.74 1.24 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.34 1.11 ;
        RECT 0.32 0.67 0.4 1.06 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.61 0.14 1.11 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OR3X4

MACRO DFFRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRXL 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 0.495 0.885 1.22 ;
        RECT 0.825 0.98 0.94 1.11 ;
        RECT 0.94 0.435 1 0.555 ;
        RECT 0.825 0.495 1 0.555 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.29 0.73 ;
        RECT 0.21 0.54 0.29 1.02 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.785 0.72 2.125 0.96 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.815 1.315 1.265 ;
        RECT 1.235 0.815 1.365 0.895 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.435 0.625 4.655 0.815 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END DFFRXL

MACRO FILL16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL16 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END FILL16

MACRO XOR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3XL 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.925 0.665 3.295 0.725 ;
        RECT 3.235 0.665 3.295 0.935 ;
        RECT 3.235 0.815 3.365 0.935 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.64 0.515 1.085 ;
        RECT 0.435 1.005 0.57 1.085 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.175 0.92 ;
        RECT 0.095 0.65 0.175 1.115 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.24 0.57 4.365 0.705 ;
        RECT 4.235 0.625 4.365 0.705 ;
        RECT 4.305 0.57 4.365 1.1 ;
        RECT 4.24 1.04 4.365 1.1 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
END XOR3XL

MACRO CLKBUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX6 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.57 1.54 1.07 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.35 0.13 1.37 ;
        RECT 0.06 0.79 0.14 0.975 ;
        RECT 0.48 0.35 0.54 0.655 ;
        RECT 0.48 0.915 0.54 1.37 ;
        RECT 0.06 0.915 0.95 0.975 ;
        RECT 0.89 0.35 0.95 0.655 ;
        RECT 0.06 0.595 0.95 0.655 ;
        RECT 0.89 0.915 0.95 1.37 ;
    END
  END Y
END CLKBUFX6

MACRO AOI222XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222XL 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 0.24 0.9 0.36 ;
        RECT 1.585 1.01 1.645 1.195 ;
        RECT 0.84 0.27 1.92 0.33 ;
        RECT 1.86 0.27 1.92 1.07 ;
        RECT 1.585 1.01 1.92 1.07 ;
        RECT 1.86 0.41 1.94 0.54 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 0.575 1.025 0.895 ;
        RECT 0.835 0.815 1.095 0.895 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.47 1.74 0.91 ;
        RECT 1.62 0.83 1.76 0.91 ;
    END
  END C1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.215 0.615 0.335 0.895 ;
        RECT 0.035 0.815 0.335 0.895 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.195 0.745 1.34 0.825 ;
        RECT 1.26 0.6 1.34 1.035 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.43 1.52 0.91 ;
        RECT 1.44 0.43 1.54 0.73 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.46 0.555 0.895 ;
        RECT 0.435 0.815 0.58 0.895 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END AOI222XL

MACRO OR4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X6 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2 0.98 2.06 1.37 ;
        RECT 2.09 0.275 2.15 0.585 ;
        RECT 2 0.98 2.74 1.04 ;
        RECT 2.41 0.98 2.47 1.37 ;
        RECT 2.5 0.275 2.56 0.585 ;
        RECT 2.66 0.525 2.72 1.11 ;
        RECT 2.41 0.98 2.74 1.11 ;
        RECT 2.41 1.05 2.88 1.11 ;
        RECT 2.82 1.05 2.88 1.37 ;
        RECT 2.91 0.275 2.97 0.585 ;
        RECT 2.09 0.525 2.97 0.585 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 0.89 0.36 1.23 ;
        RECT 1.66 0.805 1.72 1.23 ;
        RECT 0.3 1.17 1.72 1.23 ;
        RECT 1.66 0.98 1.74 1.11 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 1.07 ;
        RECT 0.46 0.92 0.58 1.07 ;
        RECT 1.5 0.89 1.56 1.07 ;
        RECT 0.46 1.01 1.56 1.07 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.625 1.365 0.705 ;
        RECT 1.305 0.625 1.365 0.91 ;
        RECT 0.68 0.85 1.365 0.91 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 0.625 0.965 0.75 ;
        RECT 0.68 0.67 1.135 0.75 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END OR4X6

MACRO ACHCONX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ACHCONX2 0 0 ;
  SIZE 7.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.03 0.815 6.09 1.13 ;
        RECT 5.515 1.07 6.09 1.13 ;
        RECT 6.115 0.325 6.175 0.895 ;
        RECT 6.03 0.815 6.175 0.895 ;
        RECT 6.03 1.015 6.545 1.075 ;
        RECT 5.385 0.325 6.63 0.385 ;
    END
  END CON
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.035 0.675 0.205 1.085 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.58 0.695 1.76 0.925 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.805 0.775 7.265 0.895 ;
    END
  END CI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.4 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.4 1.71 ;
    END
  END VDD
END ACHCONX2

MACRO OAI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.71 1.2 0.77 1.48 ;
        RECT 0.915 0.37 0.975 0.49 ;
        RECT 0.915 0.43 1.12 0.49 ;
        RECT 1.06 0.43 1.12 1.26 ;
        RECT 1.06 0.98 1.14 1.26 ;
        RECT 0.71 1.2 1.14 1.26 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.54 0.88 ;
        RECT 0.46 0.6 0.76 0.68 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 1.1 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OAI21X1

MACRO DLY3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY3X4 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.58 0.61 1.66 1.02 ;
        RECT 1.66 0.6 1.74 0.73 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.44 0.475 2.56 0.535 ;
        RECT 2.46 0.475 2.56 0.73 ;
        RECT 2.54 0.6 2.6 1.29 ;
        RECT 2.91 0.475 3.01 0.66 ;
        RECT 2.46 0.6 3.01 0.66 ;
        RECT 2.95 0.475 3.01 1.29 ;
        RECT 2.91 0.475 3.03 0.535 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.2 0.06 ;
    END
  END VSS
END DLY3X4

MACRO TLATNSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.985 0.51 4.065 0.67 ;
        RECT 4.06 0.59 4.14 1.04 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 0.9 3.115 1.04 ;
        RECT 3.06 0.51 3.14 0.98 ;
    END
  END QN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.63 4.34 1.04 ;
        RECT 4.26 0.735 4.43 1.04 ;
    END
  END GN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.75 2.74 1.25 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.49 0.79 1.94 0.87 ;
        RECT 1.86 0.79 1.94 0.92 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.755 0.61 1.025 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END TLATNSRX2

MACRO AND3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.405 1.14 1.385 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.72 0.76 0.8 1.06 ;
        RECT 0.72 0.98 0.94 1.06 ;
        RECT 0.86 0.98 0.94 1.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.98 ;
        RECT 0.38 0.6 0.46 0.91 ;
        RECT 0.26 0.79 0.46 0.91 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 1.1 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END AND3XL

MACRO DFFSXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSXL 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.49 0.94 1.02 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.305 0.73 ;
        RECT 0.225 0.54 0.305 1.02 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.66 0.46 4.74 0.96 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.46 4.54 0.96 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.73 0.815 2.185 0.895 ;
        RECT 2.035 0.815 2.185 0.94 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END DFFSXL

MACRO NAND4BBXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBXL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.69 1.23 0.75 1.385 ;
        RECT 0.555 0.36 1.175 0.42 ;
        RECT 1.06 0.98 1.175 1.29 ;
        RECT 0.69 1.23 1.175 1.29 ;
        RECT 1.115 0.36 1.175 1.385 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.815 0.7 1.13 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 0.84 0.88 1.13 ;
        RECT 0.86 0.69 0.94 0.92 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.275 0.815 1.565 0.895 ;
        RECT 1.415 0.815 1.565 1.105 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.5 0.14 0.745 ;
        RECT 0.095 0.625 0.175 0.965 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END NAND4BBXL

MACRO CLKBUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX16 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.585 0.29 0.965 ;
        RECT 0.275 0.525 0.335 0.645 ;
        RECT 0.26 0.905 0.335 1.345 ;
        RECT 0.26 0.905 0.34 1.11 ;
        RECT 0.685 0.905 0.745 1.345 ;
        RECT 0.655 0.57 0.775 0.645 ;
        RECT 1.095 0.905 1.155 1.345 ;
        RECT 1.065 0.57 1.185 0.645 ;
        RECT 1.505 0.905 1.565 1.345 ;
        RECT 1.475 0.57 1.595 0.645 ;
        RECT 1.915 0.905 1.975 1.345 ;
        RECT 1.885 0.57 2.005 0.645 ;
        RECT 2.325 0.905 2.385 1.345 ;
        RECT 2.295 0.57 2.415 0.645 ;
        RECT 0.23 0.905 2.795 0.965 ;
        RECT 0.23 0.585 2.735 0.645 ;
        RECT 2.735 0.905 2.795 1.345 ;
        RECT 2.69 0.57 2.825 0.63 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.815 3.76 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END CLKBUFX16

MACRO OAI221X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.79 1.2 0.85 1.48 ;
        RECT 0.79 1.2 1.365 1.26 ;
        RECT 1.305 1.09 1.365 1.49 ;
        RECT 1.26 1.2 1.365 1.49 ;
        RECT 1.44 0.39 1.5 1.15 ;
        RECT 1.305 1.09 1.5 1.15 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 1.1 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.6 1.14 1.1 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.47 1.34 0.97 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END OAI221X1

MACRO AND4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 0.26 1.235 0.38 ;
        RECT 1.175 0.32 1.34 0.38 ;
        RECT 1.26 0.32 1.34 0.54 ;
        RECT 1.27 0.32 1.34 1.245 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.86 1.08 1.25 ;
        RECT 1.06 1.17 1.14 1.3 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.64 0.72 1.12 ;
        RECT 0.64 0.64 0.74 0.92 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.64 0.52 1.12 ;
        RECT 0.44 0.64 0.54 0.92 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 0.64 0.34 1.1 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END AND4XL

MACRO OAI31X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.73 1.2 0.79 1.48 ;
        RECT 1.06 0.37 1.14 0.54 ;
        RECT 1.08 0.37 1.14 1.26 ;
        RECT 0.73 1.2 1.14 1.26 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.17 0.53 0.25 0.87 ;
        RECT 0.06 0.79 0.25 0.87 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 1.1 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 1.1 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OAI31X1

MACRO OA21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.6 1.14 1.455 ;
        RECT 1.08 0.57 1.3 0.63 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.56 0.14 1.06 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.59 0.54 1.09 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.22 0.74 0.72 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END OA21X1

MACRO DLY4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY4X4 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.86 0.98 5.94 1.235 ;
        RECT 5.89 0.765 5.97 1.06 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.49 0.72 0.99 ;
        RECT 0.57 0.93 0.72 0.99 ;
        RECT 0.66 0.6 0.74 0.73 ;
        RECT 0.66 0.67 1.13 0.73 ;
        RECT 1.07 0.49 1.13 0.99 ;
        RECT 1.04 0.93 1.16 0.99 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.2 0.06 ;
    END
  END VSS
END DLY4X4

MACRO CLKXOR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X8 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 0.435 0.315 0.555 ;
        RECT 0.26 0.495 0.32 1.36 ;
        RECT 0.26 0.495 0.34 0.73 ;
        RECT 0.67 0.915 0.73 1.36 ;
        RECT 0.635 0.48 0.755 0.555 ;
        RECT 1.08 0.915 1.14 1.36 ;
        RECT 1.045 0.48 1.165 0.555 ;
        RECT 0.255 0.495 1.485 0.555 ;
        RECT 0.26 0.915 1.55 0.975 ;
        RECT 1.49 0.915 1.55 1.36 ;
        RECT 1.44 0.48 1.575 0.54 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.72 0.61 3.14 0.69 ;
        RECT 3.06 0.61 3.14 0.92 ;
        RECT 3.06 0.79 3.18 0.87 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.625 2.03 0.745 ;
        RECT 1.95 0.625 2.03 1.01 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END CLKXOR2X8

MACRO OR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X8 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.225 1 1.285 1.445 ;
        RECT 1.27 0.57 1.39 0.63 ;
        RECT 1.635 1 1.695 1.445 ;
        RECT 1.68 0.57 1.8 0.645 ;
        RECT 2.045 1 2.105 1.445 ;
        RECT 2.12 0.525 2.18 0.645 ;
        RECT 2.26 0.585 2.32 1.06 ;
        RECT 2.26 0.585 2.34 0.73 ;
        RECT 1.225 1 2.515 1.06 ;
        RECT 2.455 1 2.515 1.445 ;
        RECT 1.345 0.585 2.53 0.645 ;
        RECT 2.485 0.57 2.62 0.63 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.925 0.54 1.3 ;
        RECT 0.46 0.925 0.665 1.005 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.36 0.92 ;
        RECT 0.28 0.745 0.965 0.825 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END OR2X8

MACRO DFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFXL 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.56 0.94 1.3 ;
        RECT 0.92 0.52 1 0.64 ;
        RECT 0.86 0.995 1.055 1.115 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.54 0.27 0.73 ;
        RECT 0.19 0.54 0.27 1.02 ;
        RECT 0.06 0.54 0.35 0.66 ;
        RECT 0.27 0.94 0.35 1.06 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.93 0.845 4.14 1.185 ;
        RECT 3.93 0.845 4.17 1.085 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.62 1.38 0.79 ;
        RECT 1.3 0.62 1.38 0.895 ;
        RECT 1.3 0.815 1.565 0.895 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END DFFXL

MACRO OAI2BB2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X4 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.705 1.11 1.765 1.23 ;
        RECT 1.705 1.11 2.735 1.17 ;
        RECT 2.425 1.11 2.485 1.335 ;
        RECT 2.425 1.11 2.735 1.275 ;
        RECT 2.905 0.465 2.965 1.275 ;
        RECT 2.835 1.195 2.965 1.275 ;
        RECT 3.115 0.445 3.235 0.525 ;
        RECT 2.425 1.215 3.525 1.275 ;
        RECT 3.555 0.305 3.615 0.525 ;
        RECT 2.905 0.465 3.615 0.525 ;
        RECT 3.555 0.305 3.675 0.365 ;
        RECT 4.11 0.285 4.23 0.365 ;
        RECT 3.465 1.155 4.45 1.215 ;
        RECT 3.625 0.285 4.6 0.345 ;
        RECT 4.55 0.305 4.67 0.365 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.285 0.625 3.365 0.745 ;
        RECT 3.085 0.625 3.545 0.705 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.125 0.845 3.365 1.085 ;
        RECT 3.065 0.845 4.535 0.905 ;
        RECT 4.475 0.835 4.685 0.895 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.685 0.54 1.185 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.685 0.34 1.185 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END OAI2BB2X4

MACRO EDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFX1 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.6 5.34 0.73 ;
        RECT 5.28 0.54 5.34 1.29 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.54 4.54 1.29 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.175 0.695 3.295 0.755 ;
        RECT 3.235 0.695 3.295 1.515 ;
        RECT 2.965 1.455 3.295 1.515 ;
        RECT 3.235 1.08 4.12 1.14 ;
        RECT 4.06 0.975 4.14 1.11 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.555 0.805 3.765 0.98 ;
        RECT 3.555 0.805 3.96 0.885 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 0.77 0.38 1.06 ;
        RECT 0.3 0.98 0.54 1.06 ;
        RECT 0.46 0.98 0.54 1.11 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END EDFFX1

MACRO HOLDX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HOLDX1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 0.74 0.4 0.98 ;
        RECT 0.86 0.79 0.94 0.98 ;
        RECT 0.34 0.92 0.94 0.98 ;
        RECT 0.87 0.54 0.94 1.02 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END HOLDX1

MACRO TLATNTSCAX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX8 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.96 3.74 1.11 ;
        RECT 3.68 0.515 3.74 1.405 ;
        RECT 4.09 0.96 4.15 1.405 ;
        RECT 4.06 0.545 4.18 0.605 ;
        RECT 4.5 0.96 4.56 1.405 ;
        RECT 4.47 0.545 4.59 0.62 ;
        RECT 4.135 0.56 4.97 0.62 ;
        RECT 3.66 0.96 4.97 1.02 ;
        RECT 4.91 0.5 4.97 1.405 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.74 0.73 ;
        RECT 0.675 0.6 0.755 0.935 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 0.45 0.525 0.935 ;
        RECT 0.445 0.45 0.54 0.73 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.065 0.465 0.185 0.895 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.2 0.06 ;
    END
  END VSS
END TLATNTSCAX8

MACRO ANTENNA
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ANTENNA 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.6 0.06 ;
    END
  END VSS
  PIN A
    ANTENNADIFFAREA 1.7285  LAYER Metal1 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.39 0.34 1.27 ;
    END
  END A
END ANTENNA

#MACRO ANTENNA
#  CLASS CORE ;
#  ORIGIN 0 0 ;
#  FOREIGN ANTENNA 0 0 ;
#  SIZE 0.6 BY 1.71 ;
#  SYMMETRY X Y ;
#  SITE CoreSite ;
#  PIN VDD
#    DIRECTION INOUT ;
#    USE POWER ;
#    SHAPE ABUTMENT ;
#    NETEXPR "VDD VDD!" ;
#    PORT
#      LAYER Metal1 ;
#        RECT 0.00 1.65 0.6 1.71 ;
#    END
#  END VDD
#  PIN VSS
#    DIRECTION INOUT ;
#    USE GROUND ;
#    SHAPE ABUTMENT ;
#    NETEXPR "VSS VSS!" ;
#    PORT
#      LAYER Metal1 ;
#        RECT 0.00 0.00 0.6 0.06 ;
#    END
#  END VSS
#  PIN A
#    DIRECTION INPUT ;
#    USE SIGNAL ;
#    PORT
#      LAYER Metal1 ;
#        RECT 0.26 0.39 0.34 1.27 ;
#    END
#  END A
#END ANTENNA

MACRO OAI2BB2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X1 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 1.195 1.805 1.275 ;
        RECT 1.745 1.195 1.805 1.315 ;
        RECT 1.995 0.38 2.055 0.5 ;
        RECT 2.04 0.44 2.1 1.255 ;
        RECT 1.435 1.195 2.1 1.255 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.465 2.34 0.905 ;
        RECT 2.2 0.755 2.34 0.905 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.595 1.94 1.095 ;
    END
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 0.815 0.71 1.105 ;
        RECT 0.625 1.005 0.915 1.105 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.815 0.525 0.895 ;
        RECT 0.445 0.815 0.525 1.105 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END OAI2BB2X1

MACRO CLKINVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX1 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.28 0.51 0.34 1.29 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.59 0.16 0.79 ;
        RECT 0.08 0.59 0.16 1.07 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.6 0.06 ;
    END
  END VSS
END CLKINVX1

MACRO SDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX2 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.36 0.92 ;
        RECT 0.3 0.54 0.36 1.335 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.195 0.5 4.255 0.88 ;
        RECT 4.44 0.5 4.56 0.67 ;
        RECT 5.025 0.815 5.165 0.875 ;
        RECT 4.195 0.5 5.145 0.56 ;
        RECT 5.085 0.5 5.145 0.895 ;
        RECT 5.035 0.815 5.165 0.895 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.845 0.66 4.925 0.975 ;
        RECT 4.66 0.785 4.925 0.975 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.5 3.74 0.73 ;
        RECT 3.66 0.645 3.935 0.73 ;
        RECT 3.855 0.645 3.935 0.805 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.94 0.54 1.115 ;
        RECT 0.635 0.89 0.815 1.02 ;
        RECT 0.46 0.94 0.815 1.02 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END SDFFHQX2

MACRO SDFFSRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX8 0 0 ;
  SIZE 9.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.4 0.6 8.46 0.88 ;
        RECT 8.4 0.6 9.34 0.66 ;
        RECT 9.26 0.6 9.34 0.73 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.835 0.76 9.16 0.96 ;
        RECT 8.78 0.82 9.16 0.96 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.06 0.445 8.14 0.945 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.635 0.625 7.96 0.705 ;
        RECT 7.88 0.625 7.96 0.88 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.79 3.14 0.92 ;
        RECT 3.12 0.815 3.18 1.015 ;
        RECT 3.12 0.955 4.12 1.015 ;
        RECT 4.06 0.955 4.12 1.365 ;
        RECT 4.86 1.135 4.92 1.365 ;
        RECT 4.06 1.305 4.92 1.365 ;
        RECT 4.86 1.135 5.3 1.195 ;
        RECT 5.24 1.135 5.3 1.34 ;
        RECT 5.24 1.28 6 1.34 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.565 0.79 2.765 0.975 ;
        RECT 2.565 0.79 2.96 0.87 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.54 0.14 1.345 ;
        RECT 0.49 0.54 0.55 1.345 ;
        RECT 0.06 0.6 0.96 0.66 ;
        RECT 0.9 0.54 0.96 1.345 ;
        RECT 0.9 0.74 1.325 0.8 ;
        RECT 1.265 0.59 1.325 0.96 ;
        RECT 1.31 0.53 1.37 0.65 ;
        RECT 1.31 0.9 1.37 1.345 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 9.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 9.6 0.06 ;
    END
  END VSS
END SDFFSRHQX8

MACRO CLKXOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.28 0.495 0.34 1.215 ;
        RECT 0.28 1.155 0.435 1.215 ;
        RECT 0.375 0.435 0.435 0.555 ;
        RECT 0.28 0.495 0.435 0.555 ;
        RECT 0.375 1.155 0.435 1.275 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.825 1.565 0.885 ;
        RECT 1.435 0.815 1.565 0.895 ;
        RECT 1.335 0.815 1.785 0.875 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 0.815 0.8 0.895 ;
        RECT 0.72 0.815 0.8 1.195 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END CLKXOR2X2

MACRO OAI221X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 1.21 0.63 1.33 ;
        RECT 1.45 1.21 1.51 1.33 ;
        RECT 2.425 1.21 2.485 1.33 ;
        RECT 3.045 1.21 3.105 1.33 ;
        RECT 3.715 1.07 3.775 1.46 ;
        RECT 3.805 0.535 3.865 0.675 ;
        RECT 0.57 1.21 4.185 1.27 ;
        RECT 4.125 1.07 4.185 1.46 ;
        RECT 4.215 0.535 4.3 0.675 ;
        RECT 3.805 0.615 4.3 0.675 ;
        RECT 4.24 0.535 4.3 1.13 ;
        RECT 4.125 1.07 4.3 1.13 ;
        RECT 4.24 0.79 4.34 0.92 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.22 0.86 0.34 0.92 ;
        RECT 0.28 0.79 0.34 1.055 ;
        RECT 1.01 0.935 1.07 1.055 ;
        RECT 1.695 0.91 1.755 1.055 ;
        RECT 0.28 0.995 1.755 1.055 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.09 0.875 2.15 1.11 ;
        RECT 2.77 0.94 2.89 1.11 ;
        RECT 3.46 0.91 3.54 1.11 ;
        RECT 2.09 1.05 3.54 1.11 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.615 0.775 0.765 0.895 ;
        RECT 0.615 0.775 1.475 0.835 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.47 0.775 3.12 0.835 ;
        RECT 3.035 0.815 3.165 0.895 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.64 0.815 4.14 0.895 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END OAI221X4

MACRO XNOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.925 0.665 3.295 0.725 ;
        RECT 3.235 0.665 3.295 0.935 ;
        RECT 3.235 0.815 3.365 0.935 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 0.605 0.49 0.75 ;
        RECT 0.46 0.67 0.54 1.055 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.15 0.92 ;
        RECT 0.07 0.615 0.15 1.105 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.235 0.435 4.365 0.515 ;
        RECT 4.305 0.435 4.365 0.99 ;
        RECT 4.24 0.93 4.365 0.99 ;
    END
  END Y
END XNOR3X1

MACRO SEDFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFXL 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.845 0.375 3.925 0.5 ;
        RECT 3.86 0.42 3.94 1.16 ;
        RECT 3.86 1.08 3.98 1.16 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.65 1.775 0.73 ;
        RECT 1.63 0.48 1.71 0.68 ;
        RECT 1.63 0.6 1.74 0.68 ;
        RECT 1.695 0.65 1.775 1.21 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.86 0.79 6.94 1.06 ;
        RECT 6.86 0.79 7.17 0.91 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 0.57 3.54 1.07 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.735 2.34 0.975 ;
        RECT 2.44 0.735 2.52 0.895 ;
        RECT 2.26 0.815 2.52 0.895 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.805 0.705 0.955 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.645 0.335 0.77 ;
        RECT 0.705 0.325 0.765 0.705 ;
        RECT 0.635 0.625 0.765 0.705 ;
        RECT 0.275 0.645 0.865 0.705 ;
        RECT 0.805 0.645 0.865 0.77 ;
        RECT 0.705 0.325 1.345 0.385 ;
        RECT 1.285 0.325 1.345 0.93 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.2 0.06 ;
    END
  END VSS
END SEDFFXL

MACRO OA22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.6 1.54 0.73 ;
        RECT 1.44 0.67 1.5 1.33 ;
        RECT 1.48 0.525 1.54 0.73 ;
        RECT 1.48 0.525 1.615 0.585 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.87 1.08 1.06 ;
        RECT 1 0.98 1.34 1.06 ;
        RECT 1.26 0.98 1.34 1.11 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.64 0.74 1.14 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OA22X1

MACRO AOI211X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.44 0.7 0.5 ;
        RECT 1.035 1.12 1.095 1.48 ;
        RECT 1.06 0.41 1.14 0.54 ;
        RECT 0.63 0.48 1.3 0.54 ;
        RECT 1.24 0.48 1.3 1.18 ;
        RECT 1.035 1.12 1.3 1.18 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.54 1.1 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.64 0.74 1.04 ;
        RECT 0.66 0.64 0.84 0.72 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 0.64 1.02 0.87 ;
        RECT 0.94 0.79 1.14 0.87 ;
        RECT 1.06 0.79 1.14 1.02 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END AOI211X1

MACRO TLATX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATX4 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.98 2.36 1.355 ;
        RECT 2.42 0.465 2.48 1.085 ;
        RECT 2.26 0.98 2.48 1.085 ;
        RECT 2.26 1.025 2.77 1.085 ;
        RECT 2.71 1.025 2.77 1.355 ;
        RECT 2.89 0.465 2.95 0.585 ;
        RECT 2.42 0.525 2.95 0.585 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.54 0.465 0.6 0.585 ;
        RECT 0.66 0.79 0.72 1.355 ;
        RECT 0.68 0.525 0.74 1.025 ;
        RECT 0.66 0.965 1.13 1.025 ;
        RECT 1.01 0.465 1.07 0.585 ;
        RECT 0.54 0.525 1.07 0.585 ;
        RECT 1.07 0.965 1.13 1.355 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.235 0.79 4.54 0.92 ;
        RECT 4.46 0.79 4.54 1.065 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.46 0.34 0.96 ;
    END
  END G
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END TLATX4

MACRO BUFX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX20 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.355 0.13 1.36 ;
        RECT 0.06 0.595 0.14 0.975 ;
        RECT 0.48 0.355 0.54 0.655 ;
        RECT 0.48 0.915 0.54 1.36 ;
        RECT 0.89 0.355 0.95 0.655 ;
        RECT 0.89 0.915 0.95 1.36 ;
        RECT 1.3 0.355 1.36 0.655 ;
        RECT 1.3 0.915 1.36 1.36 ;
        RECT 1.71 0.355 1.77 0.655 ;
        RECT 1.71 0.915 1.77 1.36 ;
        RECT 2.12 0.355 2.18 0.655 ;
        RECT 2.12 0.915 2.18 1.36 ;
        RECT 2.53 0.355 2.59 0.655 ;
        RECT 2.53 0.915 2.59 1.36 ;
        RECT 2.94 0.355 3 0.655 ;
        RECT 2.94 0.915 3 1.36 ;
        RECT 0.06 0.915 3.41 0.975 ;
        RECT 3.35 0.355 3.41 0.655 ;
        RECT 0.06 0.595 3.41 0.655 ;
        RECT 3.35 0.915 3.41 1.36 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.875 0.815 4.375 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END BUFX20

MACRO XNOR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2XL 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.2 0.73 ;
        RECT 0.12 0.6 0.2 1.1 ;
        RECT 0.215 0.485 0.295 0.68 ;
        RECT 0.06 0.6 0.295 0.68 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.27 0.815 1.77 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 1.075 ;
        RECT 0.565 0.68 0.645 0.87 ;
        RECT 0.46 0.79 0.645 0.87 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END XNOR2XL

MACRO OR4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.395 1.3 1.385 ;
        RECT 1.24 0.41 1.34 0.54 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.98 0.54 1.11 ;
        RECT 0.51 0.66 0.59 1.07 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 1.02 ;
        RECT 0.33 0.59 0.41 0.87 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.03 0.735 0.12 1.04 ;
        RECT 0.06 0.59 0.16 0.795 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.475 1.14 0.765 ;
        RECT 0.85 0.685 1.14 0.765 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END OR4X1

MACRO OAI211XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 1.25 1.14 1.31 ;
        RECT 1.04 0.295 1.1 1.31 ;
        RECT 1.06 1.19 1.14 1.38 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.8 0.34 1.3 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.65 0.54 1.15 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.655 0.745 0.92 ;
        RECT 0.665 0.655 0.745 1.15 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 1.1 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OAI211XL

MACRO BUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX4 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.42 0.29 1.04 ;
        RECT 0.275 0.36 0.335 0.48 ;
        RECT 0.26 0.98 0.335 1.37 ;
        RECT 0.26 0.98 0.34 1.11 ;
        RECT 0.23 0.98 0.76 1.04 ;
        RECT 0.23 0.42 0.72 0.48 ;
        RECT 0.7 0.98 0.76 1.37 ;
        RECT 0.67 0.4 0.79 0.46 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.78 0.94 1.15 ;
        RECT 0.95 0.74 1.03 0.86 ;
        RECT 0.86 0.78 1.03 0.86 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END BUFX4

MACRO CLKINVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX4 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 0.54 0.46 0.68 ;
        RECT 0.4 0.995 0.46 1.335 ;
        RECT 0.4 0.995 0.94 1.055 ;
        RECT 0.81 0.54 0.87 0.68 ;
        RECT 0.4 0.62 0.92 0.68 ;
        RECT 0.81 0.995 0.87 1.335 ;
        RECT 0.86 0.62 0.92 1.11 ;
        RECT 0.86 0.98 0.94 1.11 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.815 0.76 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END CLKINVX4

MACRO AOI33X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.64 0.335 2.7 0.92 ;
        RECT 2.64 0.79 2.74 0.92 ;
        RECT 2.64 0.815 3.03 0.895 ;
        RECT 2.97 0.815 3.03 1.115 ;
        RECT 2.97 0.995 3.44 1.055 ;
        RECT 3.38 0.995 3.44 1.205 ;
        RECT 3.79 1.085 3.85 1.205 ;
        RECT 4.2 1.085 4.26 1.205 ;
        RECT 0.955 0.335 4.6 0.395 ;
        RECT 4.61 1.085 4.67 1.205 ;
        RECT 3.38 1.085 5.08 1.145 ;
        RECT 5.02 1.085 5.08 1.205 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 0.845 1.29 0.905 ;
        RECT 1.23 0.845 1.29 0.985 ;
        RECT 1.23 0.925 2.095 0.985 ;
        RECT 2.035 0.815 2.125 0.935 ;
        RECT 2.035 0.815 2.165 0.895 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.435 0.815 3.6 0.895 ;
        RECT 3.54 0.815 3.6 0.985 ;
        RECT 4.28 0.835 4.34 0.985 ;
        RECT 3.54 0.925 4.34 0.985 ;
        RECT 4.28 0.835 4.57 0.895 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.07 0.655 3.76 0.715 ;
        RECT 3.7 0.655 3.76 0.825 ;
        RECT 4.12 0.675 4.18 0.825 ;
        RECT 3.7 0.765 4.18 0.825 ;
        RECT 4.12 0.675 4.73 0.735 ;
        RECT 4.67 0.675 4.73 0.835 ;
        RECT 4.67 0.775 4.95 0.835 ;
        RECT 4.86 0.775 4.94 0.92 ;
        RECT 4.86 0.775 4.95 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 0.79 0.74 0.85 ;
        RECT 0.68 0.685 0.74 0.92 ;
        RECT 0.66 0.79 0.74 0.92 ;
        RECT 0.68 0.685 1.45 0.745 ;
        RECT 1.39 0.685 1.45 0.825 ;
        RECT 1.875 0.655 1.935 0.825 ;
        RECT 1.39 0.765 1.935 0.825 ;
        RECT 1.875 0.655 2.36 0.715 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.495 0.5 0.695 ;
        RECT 1.55 0.495 1.67 0.665 ;
        RECT 0.44 0.495 2.54 0.555 ;
        RECT 2.46 0.495 2.54 0.73 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.905 0.495 2.965 0.665 ;
        RECT 2.8 0.585 2.965 0.665 ;
        RECT 3.9 0.495 4.02 0.665 ;
        RECT 2.905 0.495 5.11 0.555 ;
        RECT 5.05 0.495 5.11 0.705 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END AOI33X4

MACRO TBUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX16 0 0 ;
  SIZE 9 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.5 0.37 5.56 0.51 ;
        RECT 5.5 0.45 5.72 0.51 ;
        RECT 5.615 1.065 5.675 1.42 ;
        RECT 5.66 0.45 5.72 1.125 ;
        RECT 5.66 0.79 5.74 1.09 ;
        RECT 5.91 0.37 5.97 0.51 ;
        RECT 6.025 0.45 6.085 1.42 ;
        RECT 6.32 0.37 6.38 0.51 ;
        RECT 5.91 0.45 6.38 0.51 ;
        RECT 6.435 1.03 6.495 1.42 ;
        RECT 6.73 0.37 6.79 0.51 ;
        RECT 6.845 1.03 6.905 1.42 ;
        RECT 6.73 0.45 7.2 0.51 ;
        RECT 7.14 0.37 7.2 1.09 ;
        RECT 7.255 1.03 7.315 1.42 ;
        RECT 7.55 0.37 7.61 0.51 ;
        RECT 7.665 1.03 7.725 1.42 ;
        RECT 7.96 0.37 8.02 0.51 ;
        RECT 8.075 1.03 8.135 1.42 ;
        RECT 7.55 0.45 8.43 0.51 ;
        RECT 8.37 0.37 8.43 1.09 ;
        RECT 5.66 1.03 8.545 1.09 ;
        RECT 8.485 1.03 8.545 1.42 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.515 0.87 0.765 0.93 ;
        RECT 1.035 0.41 1.095 0.99 ;
        RECT 0.705 0.93 1.095 0.99 ;
        RECT 1.035 0.815 1.165 0.895 ;
        RECT 1.035 0.41 1.485 0.47 ;
        RECT 1.425 0.41 1.485 0.705 ;
        RECT 1.595 0.645 1.655 0.83 ;
        RECT 1.805 0.41 1.865 0.705 ;
        RECT 1.425 0.645 1.865 0.705 ;
        RECT 1.805 0.41 2.305 0.47 ;
        RECT 2.245 0.41 2.305 0.735 ;
        RECT 2.34 0.675 2.4 0.845 ;
        RECT 2.565 0.41 2.625 0.735 ;
        RECT 2.245 0.675 2.625 0.735 ;
        RECT 3.02 0.45 3.12 0.51 ;
        RECT 2.565 0.41 3.08 0.47 ;
        RECT 3.06 0.45 3.12 0.67 ;
        RECT 3.06 0.61 4.98 0.67 ;
        RECT 4.92 0.635 5.18 0.695 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.71 0.415 0.92 ;
        RECT 0.26 0.71 0.935 0.77 ;
        RECT 0.875 0.71 0.935 0.83 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 9 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 9 0.06 ;
    END
  END VSS
END TBUFX16

MACRO SDFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX1 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.865 0.54 0.94 0.73 ;
        RECT 0.86 0.6 0.94 0.73 ;
        RECT 0.88 0.54 0.94 1.33 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.29 0.73 ;
        RECT 0.21 0.54 0.29 1.29 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.14 0.675 5.2 0.795 ;
        RECT 5.405 0.465 5.465 0.735 ;
        RECT 5.14 0.675 5.465 0.735 ;
        RECT 5.405 0.465 6.12 0.525 ;
        RECT 6.06 0.465 6.12 0.73 ;
        RECT 6.06 0.6 6.14 0.73 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.565 0.625 5.645 0.81 ;
        RECT 5.565 0.625 5.96 0.745 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.66 0.495 4.74 0.855 ;
        RECT 4.66 0.495 4.88 0.575 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 0.735 1.965 0.96 ;
        RECT 1.8 0.735 2.155 0.815 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.2 0.75 1.28 1.11 ;
        RECT 1.06 0.98 1.28 1.11 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END SDFFRX1

MACRO DFFSRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX8 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.46 0.655 7.54 1.155 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.765 0.625 6.885 0.865 ;
        RECT 6.835 0.495 6.975 0.705 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.79 3.14 0.92 ;
        RECT 3.08 0.79 3.14 1.265 ;
        RECT 3.42 1.125 3.48 1.265 ;
        RECT 3.08 1.205 3.48 1.265 ;
        RECT 3.42 1.125 3.96 1.185 ;
        RECT 3.9 1.125 3.96 1.345 ;
        RECT 4.9 1.22 4.96 1.345 ;
        RECT 3.9 1.285 4.96 1.345 ;
        RECT 4.9 1.22 5.34 1.28 ;
        RECT 5.28 1.22 5.34 1.44 ;
        RECT 5.28 1.38 5.59 1.44 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.6 2.74 1.1 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.54 0.14 1.345 ;
        RECT 0.49 0.54 0.55 1.345 ;
        RECT 0.06 0.645 0.96 0.705 ;
        RECT 0.9 0.54 0.96 1.345 ;
        RECT 0.9 0.74 1.325 0.8 ;
        RECT 1.265 0.59 1.325 0.96 ;
        RECT 1.31 0.53 1.37 0.65 ;
        RECT 1.31 0.9 1.37 1.345 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.8 0.06 ;
    END
  END VSS
END DFFSRHQX8

MACRO AOI222X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.79 1.34 0.92 ;
        RECT 1.28 0.45 1.34 1.065 ;
        RECT 1.28 1.005 2.5 1.065 ;
        RECT 2.44 1.005 2.5 1.155 ;
        RECT 0.705 0.45 2.675 0.51 ;
        RECT 2.44 1.02 2.91 1.08 ;
        RECT 2.85 1.015 2.91 1.135 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.815 2.135 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.79 0.835 0.92 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.555 0.79 2.725 0.92 ;
        RECT 2.555 0.815 2.74 0.895 ;
    END
  END C1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.56 0.74 ;
        RECT 0.505 0.61 0.95 0.69 ;
        RECT 0.865 0.635 1.06 0.715 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.625 1.965 0.715 ;
        RECT 1.505 0.635 2.135 0.715 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.625 2.4 0.715 ;
        RECT 2.235 0.625 2.9 0.685 ;
        RECT 2.84 0.68 3.015 0.74 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END AOI222X2

MACRO NAND2BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX1 0 0 ;
  SIZE 1.00 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.005 0.15 1.085 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.59 0.805 0.770 0.965 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.62 0.165 0.705 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.80 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.80 0.06 ;
    END
  END VSS
END NAND2BX1

MACRO AOI211X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.76 0.445 0.88 0.505 ;
        RECT 1.38 0.445 1.5 0.525 ;
        RECT 1.835 0.625 1.965 0.705 ;
        RECT 1.905 0.465 1.965 1.055 ;
        RECT 1.935 0.445 2.055 0.525 ;
        RECT 2.415 0.445 2.535 0.525 ;
        RECT 2.855 0.445 2.975 0.525 ;
        RECT 1.905 0.995 3.045 1.055 ;
        RECT 2.985 0.995 3.045 1.275 ;
        RECT 0.83 0.465 3.345 0.525 ;
        RECT 2.985 1.045 3.455 1.105 ;
        RECT 3.295 0.445 3.415 0.505 ;
        RECT 3.395 1.045 3.455 1.275 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.815 1.425 0.895 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.065 0.815 2.565 0.895 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.985 0.625 3.365 0.705 ;
        RECT 3.285 0.625 3.365 0.825 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.365 0.705 ;
        RECT 0.23 0.645 1.735 0.705 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END AOI211X4

MACRO BMXIX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BMXIX4 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.53 0.13 1.65 0.19 ;
        RECT 1.59 0.19 1.875 0.25 ;
        RECT 1.815 0.19 1.875 0.855 ;
        RECT 1.815 0.625 1.965 0.855 ;
        RECT 2.345 0.735 2.405 0.855 ;
        RECT 1.815 0.795 2.405 0.855 ;
    END
  END M1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.45 1.34 0.95 ;
    END
  END A
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 0.76 0.72 0.82 ;
        RECT 0.66 0.76 0.72 1.27 ;
        RECT 0.66 0.98 0.74 1.27 ;
        RECT 0.66 1.21 1.12 1.27 ;
        RECT 1.06 1.21 1.12 1.335 ;
        RECT 1.06 1.275 2.085 1.335 ;
    END
  END S
  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.765 0.295 1.275 ;
        RECT 0.235 1.195 0.365 1.275 ;
        RECT 0.235 1.215 0.56 1.275 ;
        RECT 0.5 1.215 0.56 1.43 ;
        RECT 0.5 1.37 0.96 1.43 ;
    END
  END M0
  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.255 0.54 4.315 1.29 ;
        RECT 4.255 0.6 4.34 0.73 ;
        RECT 4.255 0.67 4.725 0.73 ;
        RECT 4.665 0.54 4.725 1.29 ;
    END
  END PPN
  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.075 0.735 3.225 0.855 ;
        RECT 3.165 0.735 3.225 1.445 ;
        RECT 3.165 1.385 3.565 1.445 ;
        RECT 3.435 1.385 3.565 1.465 ;
    END
  END X2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END BMXIX4

MACRO MX4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4XL 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.45 0.14 1.02 ;
        RECT 0.06 0.79 0.16 1.02 ;
        RECT 0.12 0.41 0.2 0.53 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.33 1.43 2.64 1.49 ;
        RECT 3.445 0.825 3.965 0.885 ;
        RECT 2.58 1.38 3.565 1.44 ;
        RECT 3.505 0.825 3.565 1.44 ;
        RECT 3.8 0.815 3.965 0.895 ;
        RECT 3.505 0.825 3.965 0.895 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.465 0.625 3.965 0.705 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.72 0.785 2.965 0.895 ;
        RECT 2.885 0.785 2.965 1.12 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.5 0.79 2.62 0.87 ;
        RECT 2.54 0.79 2.62 1.085 ;
        RECT 2.54 1.005 2.785 1.085 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.67 1.94 1.17 ;
    END
  END D
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.46 0.62 0.54 0.87 ;
        RECT 0.26 0.79 0.54 0.87 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.2 0.06 ;
    END
  END VSS
END MX4XL

MACRO TLATX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATX2 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.6 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.6 1.71 ;
    END
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.735 0.565 1.085 ;
        RECT 0.36 0.735 0.59 0.815 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.815 2.015 1.085 ;
    END
  END G
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.41 2.32 1.305 ;
        RECT 2.26 0.41 2.34 0.54 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.46 3.34 1.305 ;
    END
  END Q
END TLATX2

MACRO TBUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX8 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.25 0.99 3.31 1.29 ;
        RECT 3.3 0.45 3.36 0.64 ;
        RECT 3.3 0.58 3.52 0.64 ;
        RECT 3.46 0.58 3.52 1.05 ;
        RECT 3.25 0.99 3.52 1.05 ;
        RECT 3.46 0.79 3.54 0.96 ;
        RECT 3.66 0.9 3.72 1.29 ;
        RECT 3.71 0.45 3.77 0.59 ;
        RECT 4.07 0.9 4.13 1.29 ;
        RECT 4.12 0.45 4.18 0.59 ;
        RECT 3.46 0.9 4.54 0.96 ;
        RECT 4.48 0.53 4.54 1.29 ;
        RECT 4.53 0.45 4.59 0.59 ;
        RECT 3.71 0.53 4.59 0.59 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.815 0.765 0.92 ;
        RECT 1.33 0.27 1.39 0.92 ;
        RECT 0.59 0.86 1.39 0.92 ;
        RECT 1.33 0.27 2.89 0.33 ;
        RECT 2.83 0.265 3.03 0.325 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.655 0.34 0.92 ;
        RECT 0.22 0.86 0.34 0.92 ;
        RECT 0.865 0.655 0.985 0.755 ;
        RECT 0.26 0.655 1.23 0.715 ;
        RECT 1.17 0.64 1.23 0.76 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END TBUFX8

MACRO NAND2BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX4 0 0 ;
  SIZE 2.00 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.065 0.545 0.145 0.625 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.385 0.925 0.465 1.005 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.855 0.785 1.935 0.930 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.00 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.00 0.06 ;
    END
  END VSS
END NAND2BX4

MACRO SDFFQXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQXL 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 1.35 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.765 0.625 3.825 0.965 ;
        RECT 3.705 0.905 3.825 0.965 ;
        RECT 3.765 0.625 4.365 0.685 ;
        RECT 4.235 0.625 4.365 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.925 0.805 4.165 0.94 ;
        RECT 3.925 0.86 4.37 0.94 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 0.815 3.445 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.34 1.225 ;
        RECT 0.33 0.795 0.41 1.06 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END SDFFQXL

MACRO AOI33X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X2 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 0.335 1.56 1.085 ;
        RECT 1.435 1.005 1.565 1.085 ;
        RECT 1.435 1.025 1.795 1.085 ;
        RECT 1.735 1.025 1.795 1.165 ;
        RECT 0.755 0.335 2.195 0.395 ;
        RECT 2.16 1.045 2.22 1.165 ;
        RECT 1.735 1.045 2.65 1.105 ;
        RECT 2.59 1.045 2.65 1.165 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.815 0.965 0.92 ;
        RECT 0.685 0.815 1.16 0.895 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.895 0.815 2.14 0.93 ;
        RECT 1.895 0.815 2.36 0.895 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 0.655 2.54 0.715 ;
        RECT 2.46 0.655 2.54 0.92 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.655 0.54 0.92 ;
        RECT 0.42 0.655 1.11 0.715 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.495 0.32 0.725 ;
        RECT 0.26 0.495 1.32 0.555 ;
        RECT 1.26 0.495 1.32 0.735 ;
        RECT 1.26 0.6 1.34 0.735 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.68 0.495 1.74 0.735 ;
        RECT 1.66 0.6 1.74 0.735 ;
        RECT 1.68 0.495 2.7 0.555 ;
        RECT 2.64 0.495 2.7 0.735 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END AOI33X2

MACRO ADDFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX1 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.8 1 3.86 1.39 ;
        RECT 3.86 0.41 3.92 1.06 ;
        RECT 3.86 0.41 3.94 0.54 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.58 0.14 0.96 ;
        RECT 0.06 0.79 0.14 0.96 ;
        RECT 0.06 0.9 0.405 0.96 ;
        RECT 0.345 0.5 0.405 0.64 ;
        RECT 0.08 0.58 0.405 0.64 ;
        RECT 0.345 0.9 0.405 1.29 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.115 0.805 1.175 0.925 ;
        RECT 1.835 0.865 1.965 1.085 ;
        RECT 1.115 0.865 2.095 0.925 ;
        RECT 2.035 0.82 3.36 0.88 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.89 0.67 1.01 0.73 ;
        RECT 0.95 0.645 1.335 0.705 ;
        RECT 1.275 0.675 1.97 0.735 ;
        RECT 1.91 0.66 3.54 0.72 ;
        RECT 3.46 0.66 3.54 0.92 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.595 0.435 1.655 0.575 ;
        RECT 1.595 0.435 1.765 0.56 ;
        RECT 1.595 0.5 3.18 0.56 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END ADDFX1

MACRO SDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX8 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.535 0.695 5.595 0.965 ;
        RECT 5.535 0.695 5.685 0.755 ;
        RECT 5.625 0.645 6.4 0.705 ;
        RECT 6.235 0.625 6.4 0.705 ;
        RECT 6.34 0.625 6.4 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.865 0.805 6.165 1.01 ;
        RECT 5.865 0.805 6.24 0.885 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.65 5.14 0.92 ;
        RECT 5.06 0.79 5.275 0.92 ;
        RECT 5.195 0.79 5.275 1.015 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.72 0.59 2.83 0.895 ;
        RECT 2.555 0.815 2.83 0.895 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.54 0.13 1.345 ;
        RECT 0.07 0.54 0.14 0.73 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.48 0.54 0.54 1.345 ;
        RECT 0.06 0.67 0.95 0.73 ;
        RECT 0.89 0.54 0.95 1.345 ;
        RECT 0.89 0.74 1.315 0.8 ;
        RECT 1.255 0.59 1.315 0.96 ;
        RECT 1.3 0.53 1.36 0.65 ;
        RECT 1.3 0.9 1.36 1.345 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END SDFFHQX8

MACRO MDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX2 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.36 0.92 ;
        RECT 0.3 0.54 0.36 1.335 ;
    END
  END Q
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.195 0.5 4.255 0.88 ;
        RECT 4.44 0.5 4.56 0.67 ;
        RECT 5.025 0.815 5.165 0.875 ;
        RECT 4.195 0.5 5.145 0.56 ;
        RECT 5.085 0.5 5.145 0.895 ;
        RECT 5.035 0.815 5.165 0.895 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.845 0.66 4.925 0.975 ;
        RECT 4.66 0.785 4.925 0.975 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.5 3.74 0.73 ;
        RECT 3.66 0.645 3.935 0.73 ;
        RECT 3.855 0.645 3.935 0.805 ;
    END
  END D0
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.94 0.54 1.115 ;
        RECT 0.635 0.89 0.815 1.02 ;
        RECT 0.46 0.94 0.815 1.02 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END MDFFHQX2

MACRO MX3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.575 0.73 ;
        RECT 0.515 0.52 0.575 1.41 ;
        RECT 0.88 0.44 0.94 0.66 ;
        RECT 0.515 1.02 0.985 1.08 ;
        RECT 0.46 0.6 0.94 0.66 ;
        RECT 0.925 0.38 0.985 0.5 ;
        RECT 0.925 1.02 0.985 1.41 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.98 0.99 3.06 1.11 ;
        RECT 3.46 0.98 3.54 1.11 ;
        RECT 2.98 1.03 3.54 1.11 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.67 3.34 0.93 ;
        RECT 3.22 0.67 3.54 0.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.46 0.485 2.54 0.985 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.485 2.34 0.985 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.76 1.34 1.19 ;
        RECT 1.26 0.76 1.41 0.84 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END MX3X4

MACRO MX2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X2 0 0 ;
  SIZE 2.0 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 0.365 1.525 0.485 ;
        RECT 1.465 1.045 1.525 1.435 ;
        RECT 1.5 0.425 1.56 1.105 ;
        RECT 1.5 0.6 1.74 0.66 ;
        RECT 1.66 0.6 1.74 0.73 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.22 0.815 1.3 1.215 ;
        RECT 1.22 0.815 1.4 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.635 0.54 1.035 ;
        RECT 0.44 0.955 0.62 1.035 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.34 1.215 ;
        RECT 0.72 0.93 0.8 1.215 ;
        RECT 0.26 1.135 0.8 1.215 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END MX2X2

MACRO NAND4BBX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 1.005 1.325 1.365 ;
        RECT 1.265 1.005 1.565 1.145 ;
        RECT 1.675 1.085 1.735 1.365 ;
        RECT 2.085 1.085 2.145 1.365 ;
        RECT 2.495 1.085 2.555 1.365 ;
        RECT 2.905 1.085 2.965 1.365 ;
        RECT 3.315 1.085 3.375 1.365 ;
        RECT 3.725 1.085 3.785 1.365 ;
        RECT 3.855 0.42 3.915 1.145 ;
        RECT 1.265 1.085 4.195 1.145 ;
        RECT 4.135 1.085 4.195 1.365 ;
        RECT 4.265 0.42 4.325 0.56 ;
        RECT 3.855 0.5 4.325 0.56 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.5 3.74 0.73 ;
        RECT 3.675 0.65 3.755 0.985 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.84 0.705 2.92 0.985 ;
        RECT 2.84 0.74 3.14 0.985 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.76 0.54 1.26 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.76 0.34 1.26 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END NAND4BBX4

MACRO BMXIX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BMXIX2 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.54 4.14 1.29 ;
    END
  END PPN
  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.525 3.74 1.025 ;
    END
  END X2
  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 0.815 2.28 0.895 ;
    END
  END M1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.165 0.88 1.315 0.96 ;
        RECT 1.235 0.655 1.44 0.895 ;
    END
  END A
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 0.995 0.565 1.085 ;
        RECT 0.435 1.005 0.565 1.085 ;
        RECT 0.505 1.035 0.63 1.095 ;
        RECT 0.57 1.035 0.63 1.44 ;
        RECT 0.57 1.38 2.005 1.44 ;
    END
  END S
  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 0.815 0.33 0.935 ;
        RECT 0.235 0.815 0.745 0.895 ;
        RECT 0.665 0.815 0.745 0.935 ;
    END
  END M0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END BMXIX2

MACRO AOI2BB1X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.45 0.14 1.105 ;
        RECT 0.43 0.37 0.49 0.51 ;
        RECT 0.08 1.045 0.695 1.105 ;
        RECT 0.635 1.045 0.695 1.43 ;
        RECT 0.84 0.37 0.9 0.51 ;
        RECT 0.08 0.45 0.9 0.51 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.705 0.54 0.92 ;
        RECT 0.36 0.705 0.96 0.785 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.45 1.14 0.73 ;
        RECT 1.12 0.6 1.2 0.89 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.565 1.54 1.065 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END AOI2BB1X2

MACRO TBUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX6 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.25 0.99 3.31 1.29 ;
        RECT 3.3 0.45 3.36 0.64 ;
        RECT 3.3 0.58 3.52 0.64 ;
        RECT 3.46 0.58 3.52 1.05 ;
        RECT 3.25 0.99 3.52 1.05 ;
        RECT 3.46 0.79 3.54 0.96 ;
        RECT 3.66 0.9 3.72 1.29 ;
        RECT 3.71 0.45 3.77 0.59 ;
        RECT 3.46 0.9 4.13 0.96 ;
        RECT 4.07 0.53 4.13 1.29 ;
        RECT 4.12 0.45 4.18 0.59 ;
        RECT 3.71 0.53 4.18 0.59 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.815 0.765 0.92 ;
        RECT 1.33 0.27 1.39 0.92 ;
        RECT 0.59 0.86 1.39 0.92 ;
        RECT 1.33 0.27 2.89 0.33 ;
        RECT 2.83 0.265 3.03 0.325 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.655 0.34 0.92 ;
        RECT 0.22 0.86 0.34 0.92 ;
        RECT 0.865 0.655 0.985 0.755 ;
        RECT 0.26 0.655 1.23 0.715 ;
        RECT 1.17 0.64 1.23 0.76 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END TBUFX6

MACRO TBUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX12 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.1 0.415 4.16 0.555 ;
        RECT 4.1 0.495 4.32 0.555 ;
        RECT 4.215 1.02 4.275 1.405 ;
        RECT 4.26 0.495 4.32 1.08 ;
        RECT 4.26 0.79 4.34 0.92 ;
        RECT 4.51 0.415 4.57 0.555 ;
        RECT 4.625 0.495 4.685 1.405 ;
        RECT 4.92 0.415 4.98 0.555 ;
        RECT 4.51 0.495 4.98 0.555 ;
        RECT 5.035 0.86 5.095 1.405 ;
        RECT 5.33 0.415 5.39 0.555 ;
        RECT 5.445 0.86 5.505 1.405 ;
        RECT 5.74 0.415 5.8 0.555 ;
        RECT 5.855 0.495 5.915 1.405 ;
        RECT 6.15 0.415 6.21 0.555 ;
        RECT 5.33 0.495 6.21 0.555 ;
        RECT 4.26 0.86 6.325 0.92 ;
        RECT 6.265 0.86 6.325 1.405 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.805 0.765 0.895 ;
        RECT 0.9 0.295 0.96 0.865 ;
        RECT 0.54 0.805 0.96 0.865 ;
        RECT 0.9 0.295 1.34 0.355 ;
        RECT 1.28 0.295 1.34 0.675 ;
        RECT 1.66 0.29 1.72 0.675 ;
        RECT 1.28 0.615 1.72 0.675 ;
        RECT 1.66 0.29 2.125 0.35 ;
        RECT 2.065 0.29 2.125 0.705 ;
        RECT 2.065 0.645 2.42 0.705 ;
        RECT 2.36 0.645 2.42 0.865 ;
        RECT 3.72 0.745 3.78 0.865 ;
        RECT 2.36 0.805 3.78 0.865 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.625 0.44 0.78 ;
        RECT 0.72 0.585 0.8 0.705 ;
        RECT 0.36 0.625 0.8 0.705 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END TBUFX12

MACRO NAND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.425 1.2 0.485 1.48 ;
        RECT 0.745 0.38 0.805 0.5 ;
        RECT 0.745 0.44 0.92 0.5 ;
        RECT 0.425 1.2 0.94 1.26 ;
        RECT 0.86 0.44 0.92 1.49 ;
        RECT 0.86 1.2 0.94 1.49 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 1.1 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.48 0.48 0.56 0.89 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END NAND3X1

MACRO DFFSRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX2 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.415 0.54 0.475 1.3 ;
        RECT 0.415 1.195 0.565 1.275 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.6 6.34 1.1 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.635 0.625 5.715 0.85 ;
        RECT 5.41 0.77 5.715 0.85 ;
        RECT 5.635 0.625 5.765 0.705 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 1.005 1.765 1.085 ;
        RECT 1.7 0.83 1.76 1.085 ;
        RECT 1.705 1.005 1.765 1.28 ;
        RECT 1.705 1.22 2.085 1.28 ;
        RECT 2.025 1.2 2.59 1.26 ;
        RECT 2.53 1.2 2.59 1.34 ;
        RECT 3.545 1.2 3.605 1.34 ;
        RECT 2.53 1.28 3.605 1.34 ;
        RECT 3.545 1.2 3.985 1.26 ;
        RECT 3.925 1.2 3.985 1.45 ;
        RECT 3.925 1.39 4.325 1.45 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.83 1.34 1.135 ;
        RECT 1.26 0.83 1.535 0.91 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END DFFSRHQX2

MACRO NAND4BBX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX1 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.85 1.2 0.91 1.48 ;
        RECT 1.26 0.98 1.34 1.26 ;
        RECT 0.85 1.2 1.34 1.26 ;
        RECT 0.615 0.305 1.345 0.365 ;
        RECT 1.28 0.98 1.34 1.48 ;
        RECT 1.285 0.305 1.345 1.085 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.485 0.625 0.565 0.905 ;
        RECT 0.435 0.815 0.565 0.905 ;
        RECT 0.485 0.625 0.735 0.705 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 0.625 0.915 1.1 ;
        RECT 0.835 0.79 0.94 1.1 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.675 0.775 1.765 0.895 ;
        RECT 1.635 0.815 1.765 0.895 ;
        RECT 1.685 0.775 1.765 1.225 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.03 0.6 0.14 0.73 ;
        RECT 0.06 0.6 0.14 1.035 ;
        RECT 0.06 0.88 0.175 1.035 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END NAND4BBX1

MACRO DFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX1 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.175 0.73 ;
        RECT 0.115 0.52 0.175 1.48 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.11 0.735 3.37 1.055 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.76 0.54 1.26 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.6 0.06 ;
    END
  END VSS
END DFFHQX1

MACRO SEDFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRXL 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.375 0.745 5.455 1.04 ;
        RECT 5.46 0.39 5.54 0.825 ;
        RECT 5.375 0.745 5.54 0.825 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 1.02 ;
        RECT 0.06 0.41 0.165 0.635 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.66 0.98 7.74 1.215 ;
        RECT 7.68 0.735 7.76 1.06 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.035 0.77 7.165 0.895 ;
        RECT 6.94 0.77 7.395 0.85 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.86 0.935 5.94 1.25 ;
        RECT 5.805 0.935 6.07 1.015 ;
    END
  END RN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.175 0.745 4.375 0.945 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.835 0.625 4.075 0.705 ;
        RECT 4.015 0.585 4.755 0.645 ;
        RECT 4.695 0.585 4.755 0.705 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.22 0.735 3.3 1.12 ;
        RECT 3.22 0.74 3.415 0.895 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8 0.06 ;
    END
  END VSS
END SEDFFTRXL

MACRO TLATNTSCAX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX6 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.35 3.92 1.37 ;
        RECT 3.86 0.76 3.94 0.92 ;
        RECT 4.27 0.35 4.33 1.37 ;
        RECT 3.86 0.76 4.74 0.82 ;
        RECT 4.635 0.6 4.695 0.82 ;
        RECT 4.68 0.35 4.74 0.66 ;
        RECT 4.68 0.76 4.74 1.37 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.74 0.95 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.45 0.54 0.95 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.48 0.2 0.895 ;
        RECT 0.035 0.815 0.2 0.895 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END TLATNTSCAX6

MACRO SDFFRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX4 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.18 0.495 6.3 0.665 ;
        RECT 6.18 0.495 6.895 0.555 ;
        RECT 6.835 0.495 6.895 0.705 ;
        RECT 6.835 0.625 6.965 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.655 0.655 6.735 0.96 ;
        RECT 6.46 0.79 6.735 0.96 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.57 0.625 5.895 0.705 ;
        RECT 5.815 0.625 5.895 0.88 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.715 0.335 1.775 0.755 ;
        RECT 1.66 0.6 1.775 0.755 ;
        RECT 2.205 0.335 2.265 0.745 ;
        RECT 1.715 0.335 3.6 0.395 ;
        RECT 3.54 0.335 3.6 0.905 ;
        RECT 3.87 0.76 3.93 0.905 ;
        RECT 3.54 0.845 3.93 0.905 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.685 0.34 1.185 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.52 0.94 0.73 ;
        RECT 0.88 0.52 0.94 1.02 ;
        RECT 0.695 0.96 0.94 1.02 ;
        RECT 0.86 0.6 1.285 0.66 ;
        RECT 1.225 0.55 1.285 1.02 ;
        RECT 1.165 0.96 1.285 1.02 ;
        RECT 1.225 0.55 1.36 0.61 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.2 0.06 ;
    END
  END VSS
END SDFFRHQX4

MACRO NAND2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2XL 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.46 0.48 0.7 0.54 ;
        RECT 0.64 0.48 0.7 1.2 ;
        RECT 0.3 1.14 0.7 1.2 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 1.02 ;
        RECT 0.18 0.64 0.26 0.92 ;
        RECT 0.06 0.79 0.26 0.92 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.395 0.64 0.54 1.04 ;
        RECT 0.36 0.79 0.54 1.04 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.8 0.06 ;
    END
  END VSS
END NAND2XL

MACRO TBUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX4 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.945 0.41 2.005 0.55 ;
        RECT 2.045 1.09 2.105 1.33 ;
        RECT 2.06 0.49 2.12 1.15 ;
        RECT 2.06 0.79 2.14 1 ;
        RECT 2.355 0.41 2.415 0.55 ;
        RECT 1.945 0.49 2.415 0.55 ;
        RECT 2.06 0.94 2.515 1 ;
        RECT 2.455 0.94 2.515 1.33 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 0.28 0.895 0.89 ;
        RECT 0.445 0.83 0.895 0.89 ;
        RECT 0.835 0.625 0.965 0.705 ;
        RECT 0.835 0.28 1.64 0.34 ;
        RECT 1.58 0.28 1.64 0.67 ;
        RECT 1.52 0.61 1.64 0.67 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 0.65 0.345 0.77 ;
        RECT 0.46 0.6 0.54 0.73 ;
        RECT 0.265 0.65 0.735 0.73 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END TBUFX4

MACRO AOI2BB2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2XL 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.87 0.655 1.95 0.935 ;
        RECT 1.87 0.815 2.17 0.895 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.625 1.61 0.705 ;
        RECT 1.53 0.625 1.61 0.835 ;
    END
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.46 0.565 0.54 ;
        RECT 0.475 0.46 0.565 0.91 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.64 0.34 1.14 ;
    END
  END A1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.08 0.465 1.14 0.73 ;
        RECT 1.06 0.6 1.14 0.73 ;
        RECT 1.08 0.465 1.77 0.525 ;
        RECT 1.71 0.465 1.77 1.095 ;
        RECT 1.71 1.035 1.83 1.095 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END AOI2BB2XL

MACRO SDFFNSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRXL 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.41 1.115 1.3 ;
        RECT 0.86 1.17 1.115 1.3 ;
        RECT 1.095 0.37 1.175 0.49 ;
        RECT 0.86 1.18 1.175 1.3 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.02 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.085 0.665 7.145 1.05 ;
        RECT 7.085 0.665 7.31 0.785 ;
        RECT 7.085 0.665 7.705 0.725 ;
        RECT 7.645 0.625 7.705 0.745 ;
        RECT 7.635 0.625 7.765 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.415 0.855 7.765 0.935 ;
        RECT 7.635 0.855 7.765 1.085 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.635 0.815 6.765 1.085 ;
        RECT 6.515 1.005 6.825 1.085 ;
    END
  END D
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.215 0.825 6.295 1.085 ;
        RECT 6.215 0.825 6.415 0.905 ;
        RECT 6.215 1.005 6.415 1.085 ;
    END
  END CKN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.825 2.32 1.11 ;
        RECT 2.28 0.98 2.34 1.235 ;
        RECT 2.28 1.175 4.41 1.235 ;
        RECT 4.35 1.175 4.41 1.365 ;
        RECT 4.35 1.305 4.805 1.365 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.75 1.565 1.12 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8 0.06 ;
    END
  END VSS
END SDFFNSRXL

MACRO ADDFHX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.605 0.435 1.765 0.55 ;
        RECT 1.605 0.49 2.27 0.55 ;
        RECT 2.21 0.55 3.38 0.61 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.88 0.655 1.975 0.715 ;
        RECT 1.915 0.71 3.78 0.77 ;
        RECT 3.66 0.71 3.74 0.92 ;
        RECT 3.66 0.71 3.78 0.79 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.87 3.56 0.895 ;
        RECT 1.135 0.815 1.815 0.875 ;
        RECT 1.755 0.87 3.56 0.93 ;
        RECT 3.5 0.87 3.56 0.99 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.6 0.14 0.98 ;
        RECT 0.08 0.92 0.405 0.98 ;
        RECT 0.345 0.52 0.405 0.66 ;
        RECT 0.06 0.6 0.405 0.66 ;
        RECT 0.345 0.92 0.405 1.29 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.1 0.54 4.16 1.29 ;
        RECT 4.1 0.6 4.34 0.73 ;
    END
  END S
END ADDFHX1

MACRO SDFFRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX1 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.175 0.73 ;
        RECT 0.095 0.45 0.175 1.41 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.58 0.645 4.64 1 ;
        RECT 4.58 0.645 5.41 0.705 ;
        RECT 5.235 0.625 5.365 0.705 ;
        RECT 5.35 0.645 5.41 0.765 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.91 0.805 5.165 1.045 ;
        RECT 4.91 0.805 5.25 0.885 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.6 4.14 0.73 ;
        RECT 4.06 0.6 4.32 0.68 ;
        RECT 4.24 0.6 4.32 0.87 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.32 0.77 1.515 0.85 ;
        RECT 1.435 0.815 1.645 1.025 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.69 0.54 1.19 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END SDFFRHQX1

MACRO CLKMX2X3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X3 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.73 0.47 1.865 0.53 ;
        RECT 1.76 0.995 1.82 1.365 ;
        RECT 1.805 0.47 1.865 1.055 ;
        RECT 1.805 0.79 1.94 0.92 ;
        RECT 1.805 0.86 2.23 0.92 ;
        RECT 2.17 0.44 2.23 0.58 ;
        RECT 1.805 0.52 2.23 0.58 ;
        RECT 2.17 0.86 2.23 1.365 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.79 1.515 1.1 ;
        RECT 1.435 0.815 1.705 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.79 0.795 0.87 ;
        RECT 0.635 0.79 0.795 1.015 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.28 0.79 0.34 1.175 ;
        RECT 0.895 0.84 0.955 1.175 ;
        RECT 0.28 1.115 0.955 1.175 ;
        RECT 0.895 0.84 1.015 0.9 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END CLKMX2X3

MACRO EDFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRX1 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 1 0.73 ;
        RECT 0.94 0.6 1 1.16 ;
        RECT 0.95 0.505 1.01 0.64 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.29 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.86 0.735 6.94 1.11 ;
        RECT 6.735 0.98 6.94 1.11 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.83 0.79 6.365 0.87 ;
        RECT 6.235 0.79 6.365 0.895 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.71 0.79 4.94 0.87 ;
        RECT 4.86 0.79 4.94 1.14 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.98 1.34 1.19 ;
        RECT 1.27 0.7 1.35 1.06 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.2 0.06 ;
    END
  END VSS
END EDFFTRX1

MACRO DFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX1 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.54 0.94 0.73 ;
        RECT 0.88 0.54 0.94 1.34 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.285 0.73 ;
        RECT 0.205 0.54 0.285 1.29 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.635 0.89 3.715 1.085 ;
        RECT 3.495 1.005 3.88 1.085 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.2 0.82 1.28 1.135 ;
        RECT 1.06 0.98 1.28 1.135 ;
        RECT 1.205 0.78 1.285 0.9 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.2 0.06 ;
    END
  END VSS
END DFFX1

MACRO MDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX8 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.535 0.695 5.595 0.965 ;
        RECT 5.535 0.695 5.685 0.755 ;
        RECT 5.625 0.645 6.4 0.705 ;
        RECT 6.235 0.625 6.4 0.705 ;
        RECT 6.34 0.625 6.4 0.745 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.865 0.805 6.165 1.01 ;
        RECT 5.865 0.805 6.24 0.885 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.65 5.14 0.92 ;
        RECT 5.06 0.79 5.275 0.92 ;
        RECT 5.195 0.79 5.275 1.015 ;
    END
  END D0
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.72 0.59 2.83 0.895 ;
        RECT 2.555 0.815 2.83 0.895 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.54 0.13 1.345 ;
        RECT 0.07 0.54 0.14 0.73 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.48 0.54 0.54 1.345 ;
        RECT 0.06 0.67 0.95 0.73 ;
        RECT 0.89 0.54 0.95 1.345 ;
        RECT 0.89 0.74 1.315 0.8 ;
        RECT 1.255 0.59 1.315 0.96 ;
        RECT 1.3 0.53 1.36 0.65 ;
        RECT 1.3 0.9 1.36 1.345 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END MDFFHQX8

MACRO CLKAND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X8 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.865 0.51 1.985 0.57 ;
        RECT 1.95 0.945 2.01 1.39 ;
        RECT 2.275 0.51 2.395 0.585 ;
        RECT 2.36 0.945 2.42 1.39 ;
        RECT 2.685 0.51 2.805 0.585 ;
        RECT 2.77 0.945 2.83 1.39 ;
        RECT 3.06 0.525 3.12 1.005 ;
        RECT 1.925 0.525 3.125 0.585 ;
        RECT 3.06 0.79 3.14 1.005 ;
        RECT 1.95 0.945 3.24 1.005 ;
        RECT 3.08 0.51 3.215 0.57 ;
        RECT 3.18 0.945 3.24 1.39 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.61 0.815 1.365 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.365 0.715 ;
        RECT 0.235 0.655 1.605 0.715 ;
        RECT 1.545 0.655 1.605 0.775 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END CLKAND2X8

MACRO CLKINVX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX20 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.355 0.335 0.66 ;
        RECT 0.275 0.92 0.335 1.36 ;
        RECT 0.685 0.355 0.745 0.66 ;
        RECT 0.685 0.92 0.745 1.36 ;
        RECT 0.275 1.08 1.155 1.14 ;
        RECT 1.095 0.355 1.155 0.66 ;
        RECT 1.095 0.92 1.155 1.36 ;
        RECT 1.505 0.355 1.565 0.66 ;
        RECT 1.505 0.92 1.565 1.36 ;
        RECT 1.915 0.355 1.975 0.66 ;
        RECT 1.915 0.92 1.975 1.36 ;
        RECT 2.325 0.355 2.385 0.66 ;
        RECT 2.325 0.92 2.385 1.36 ;
        RECT 2.735 0.355 2.795 0.66 ;
        RECT 2.735 0.92 2.795 1.36 ;
        RECT 3.145 0.355 3.205 0.66 ;
        RECT 3.145 0.92 3.205 1.36 ;
        RECT 3.3 0.6 3.36 0.98 ;
        RECT 3.46 0.79 3.54 0.98 ;
        RECT 3.555 0.355 3.615 0.66 ;
        RECT 0.275 0.6 3.615 0.66 ;
        RECT 1.095 0.92 3.7 0.98 ;
        RECT 3.64 0.905 3.7 1.36 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.76 0.565 0.895 ;
        RECT 0.32 0.76 3.105 0.82 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END CLKINVX20

MACRO OA21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 0.65 1.13 1.185 ;
        RECT 1.05 0.65 1.34 0.73 ;
        RECT 1.26 0.57 1.38 0.65 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.56 0.34 1.06 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.22 0.74 0.72 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END OA21XL

MACRO OAI211X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X2 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 1.06 0.7 1.345 ;
        RECT 1.28 0.635 1.34 1.12 ;
        RECT 1.26 0.98 1.34 1.12 ;
        RECT 1.34 1.06 1.4 1.345 ;
        RECT 0.64 1.06 1.81 1.12 ;
        RECT 1.75 1.06 1.81 1.345 ;
        RECT 1.955 0.455 2.015 0.695 ;
        RECT 1.28 0.635 2.015 0.695 ;
        RECT 1.955 0.455 2.13 0.515 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.815 0.54 1.11 ;
        RECT 0.46 0.815 0.745 0.895 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.28 0.635 0.36 0.88 ;
        RECT 0.28 0.635 0.975 0.715 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.795 1.855 0.96 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.115 0.615 2.195 0.895 ;
        RECT 2.115 0.79 2.34 0.895 ;
        RECT 2.26 0.79 2.34 0.97 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END OAI211X2

MACRO TBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX2 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.37 1.94 0.49 ;
        RECT 1.86 0.37 1.94 1.28 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.805 0.695 0.865 ;
        RECT 0.635 0.815 0.765 0.895 ;
        RECT 0.705 0.815 0.765 1.2 ;
        RECT 1.4 0.69 1.46 1.2 ;
        RECT 0.705 1.14 1.46 1.2 ;
        RECT 1.4 0.69 1.52 0.75 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.625 0.405 0.745 ;
        RECT 0.235 0.625 0.765 0.705 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END TBUFX2

MACRO DFFSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX4 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.985 0.915 7.045 1.305 ;
        RECT 7.06 0.45 7.14 0.975 ;
        RECT 6.985 0.915 7.485 0.975 ;
        RECT 7.425 0.915 7.485 1.305 ;
        RECT 6.955 0.45 7.545 0.51 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.06 0.6 6.12 1.305 ;
        RECT 6.08 0.44 6.14 0.975 ;
        RECT 6.06 0.915 6.555 0.975 ;
        RECT 6.495 0.915 6.555 1.305 ;
        RECT 6.015 0.44 6.605 0.5 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.235 0.63 3.51 0.895 ;
        RECT 3.195 0.815 3.51 0.895 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.835 0.63 3.095 0.895 ;
        RECT 2.78 0.815 3.095 0.895 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.825 0.765 1.085 ;
        RECT 0.445 1.005 0.765 1.085 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.63 0.34 1.13 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.2 0.06 ;
    END
  END VSS
END DFFSRX4

MACRO ADDHX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX1 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.81 0.51 2.89 0.63 ;
        RECT 2.81 0.89 2.89 1.29 ;
        RECT 2.86 0.55 2.94 0.97 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.235 0.73 ;
        RECT 0.175 0.415 0.235 1.47 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 0.625 1.05 0.705 ;
        RECT 0.685 0.625 1.05 0.82 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 0.465 0.565 0.705 ;
        RECT 0.435 0.625 0.565 0.705 ;
        RECT 0.6 0.285 0.66 0.525 ;
        RECT 0.445 0.465 0.66 0.525 ;
        RECT 0.6 0.285 1.53 0.345 ;
        RECT 1.47 0.285 1.53 0.435 ;
        RECT 1.47 0.375 1.91 0.435 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END ADDHX1

MACRO EDFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFXL 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.47 0.415 5.54 1.145 ;
        RECT 5.46 0.79 5.54 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.42 0.57 4.54 0.65 ;
        RECT 4.45 0.75 4.53 1.02 ;
        RECT 4.46 0.57 4.54 0.8 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.435 0.705 3.495 1.465 ;
        RECT 3.17 1.405 3.495 1.465 ;
        RECT 4.04 0.86 4.1 1.32 ;
        RECT 3.435 1.26 4.1 1.32 ;
        RECT 4.06 0.79 4.14 0.92 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.765 0.755 3.94 1.16 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.765 0.34 1.265 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END EDFFXL

MACRO OAI21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 1.2 0.7 1.385 ;
        RECT 0.755 0.38 0.815 0.5 ;
        RECT 0.755 0.44 0.92 0.5 ;
        RECT 0.86 0.44 0.92 1.26 ;
        RECT 0.86 0.98 0.94 1.26 ;
        RECT 0.64 1.2 0.94 1.26 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.76 0.14 1.26 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.8 0.54 1.3 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 1.1 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END OAI21XL

MACRO MX2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X8 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2 0.53 2.12 0.59 ;
        RECT 2.035 0.99 2.095 1.435 ;
        RECT 2.06 0.53 2.12 1.11 ;
        RECT 2.06 0.98 2.14 1.11 ;
        RECT 2.445 0.99 2.505 1.435 ;
        RECT 2.415 0.54 2.535 0.6 ;
        RECT 2.855 0.99 2.915 1.435 ;
        RECT 2.825 0.54 2.945 0.615 ;
        RECT 2.49 0.555 3.325 0.615 ;
        RECT 2.035 0.99 3.325 1.05 ;
        RECT 3.265 0.495 3.325 1.435 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 0.85 1.74 0.93 ;
        RECT 1.66 0.85 1.74 1.19 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.715 0.8 1.085 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.955 0.535 1.11 ;
        RECT 0.475 0.955 0.535 1.245 ;
        RECT 0.9 0.865 0.96 1.245 ;
        RECT 0.475 1.185 0.96 1.245 ;
        RECT 0.9 0.865 1.02 0.925 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END MX2X8

MACRO CLKMX2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X6 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.61 0.295 1.67 0.415 ;
        RECT 1.635 0.83 1.695 1.395 ;
        RECT 1.655 0.355 1.715 0.88 ;
        RECT 1.655 0.6 1.74 0.88 ;
        RECT 2.02 0.235 2.08 0.66 ;
        RECT 2.045 0.6 2.105 1.395 ;
        RECT 1.655 0.6 2.47 0.66 ;
        RECT 2.41 0.485 2.47 0.985 ;
        RECT 2.43 0.235 2.49 0.545 ;
        RECT 2.455 0.925 2.515 1.395 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.675 1.34 1.175 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.615 0.66 0.995 ;
        RECT 0.46 0.79 0.66 0.995 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.915 0.36 1.11 ;
        RECT 0.76 0.915 0.84 1.175 ;
        RECT 0.28 1.095 0.84 1.175 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END CLKMX2X6

MACRO EDFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRX4 0 0 ;
  SIZE 8.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.79 7.34 0.92 ;
        RECT 7.28 0.435 7.34 0.99 ;
        RECT 7.28 0.435 7.345 0.575 ;
        RECT 7.695 0.435 7.755 0.575 ;
        RECT 7.28 0.515 7.755 0.575 ;
        RECT 7.28 0.93 7.89 0.99 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.465 0.435 6.525 0.575 ;
        RECT 6.66 0.515 6.72 0.99 ;
        RECT 6.66 0.79 6.74 0.99 ;
        RECT 6.875 0.435 6.935 0.575 ;
        RECT 6.465 0.515 6.935 0.575 ;
        RECT 6.36 0.93 6.95 0.99 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.435 0.63 5.655 0.96 ;
        RECT 5.435 0.815 5.66 0.96 ;
        RECT 5.41 0.88 5.66 0.96 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 0.815 2.965 0.965 ;
        RECT 2.68 0.815 3.11 0.895 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.805 0.765 1.275 ;
        RECT 0.635 1.195 0.765 1.275 ;
        RECT 1.305 0.86 1.365 1.275 ;
        RECT 0.635 1.215 1.365 1.275 ;
        RECT 1.305 0.86 1.45 0.92 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.97 ;
        RECT 0.525 0.735 0.605 0.92 ;
        RECT 0.26 0.79 0.605 0.92 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.4 0.06 ;
    END
  END VSS
END EDFFTRX4

MACRO NOR2BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.45 0.14 1.27 ;
        RECT 0.08 1.21 0.31 1.27 ;
        RECT 0.25 1.21 0.31 1.33 ;
        RECT 0.31 0.43 0.415 0.49 ;
        RECT 0.08 0.45 0.37 0.51 ;
        RECT 0.355 0.37 0.415 0.49 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.815 0.765 0.895 ;
        RECT 0.685 0.75 0.765 1.005 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END NOR2BX1

MACRO SDFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX1 0 0 ;
  SIZE 7.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 0.73 ;
        RECT 0.88 0.44 0.94 0.89 ;
        RECT 0.895 0.365 0.955 0.485 ;
        RECT 0.895 0.83 0.955 1.43 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.32 0.73 ;
        RECT 0.24 0.54 0.32 1.29 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.355 0.655 6.415 1 ;
        RECT 6.675 0.595 6.735 0.715 ;
        RECT 6.835 0.625 7.14 0.715 ;
        RECT 6.355 0.655 7.14 0.715 ;
        RECT 7.08 0.625 7.14 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.635 0.815 6.98 0.93 ;
        RECT 6.515 0.85 6.98 0.93 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.595 0.815 6.095 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.605 1.005 5.765 1.085 ;
        RECT 5.685 0.995 6.095 1.075 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.995 0.815 2.165 0.875 ;
        RECT 2.035 0.815 2.165 0.985 ;
        RECT 2.035 0.925 3.045 0.985 ;
        RECT 2.985 0.925 3.045 1.215 ;
        RECT 2.985 1.155 3.945 1.215 ;
        RECT 3.885 1.155 3.945 1.375 ;
        RECT 3.885 1.315 4.4 1.375 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.71 1.34 1.21 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.4 0.06 ;
    END
  END VSS
END SDFFSRX1

MACRO CLKAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X2 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.3 0.765 0.42 ;
        RECT 0.705 0.82 0.765 1.34 ;
        RECT 0.705 0.36 0.86 0.42 ;
        RECT 0.8 0.36 0.86 0.88 ;
        RECT 0.705 0.82 0.86 0.88 ;
        RECT 0.8 0.6 0.94 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 0.68 0.485 1.06 ;
        RECT 0.46 0.98 0.54 1.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 1.29 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END CLKAND2X2

MACRO OAI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.79 0.74 0.92 ;
        RECT 0.68 0.75 0.74 1.46 ;
        RECT 0.68 0.75 0.895 0.81 ;
        RECT 0.835 0.58 0.895 0.81 ;
        RECT 0.905 0.52 0.965 0.64 ;
        RECT 0.835 0.58 0.965 0.64 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.75 0.56 1.23 ;
        RECT 0.46 0.9 0.56 1.23 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.12 0.75 0.34 0.83 ;
        RECT 0.26 0.75 0.34 1.11 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.74 1.14 1.24 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 0.91 0.92 1.23 ;
        RECT 0.86 1.17 0.94 1.39 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END OAI22X1

MACRO DFFSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX2 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.57 7.34 1.11 ;
        RECT 7.285 0.915 7.365 1.305 ;
        RECT 7.26 0.57 7.455 0.65 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.86 0.98 6.96 1.11 ;
        RECT 6.88 0.54 6.96 1.305 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.54 0.705 6.62 1.085 ;
        RECT 6.42 1.005 6.62 1.085 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.815 1.995 1.065 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 0.815 0.965 1.03 ;
        RECT 0.655 0.95 1.02 1.03 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.06 0.46 0.235 0.54 ;
        RECT 0.155 0.46 0.235 0.815 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8 0.06 ;
    END
  END VSS
END DFFSRX2

MACRO OAI32X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.79 0.94 0.92 ;
        RECT 0.88 0.65 0.94 1.36 ;
        RECT 1.2 0.44 1.26 0.71 ;
        RECT 0.88 0.65 1.26 0.71 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.52 0.34 1.02 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.8 0.54 1.3 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.81 1.14 1.31 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.98 0.74 1.13 ;
        RECT 0.68 0.65 0.76 1.04 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.36 0.52 1.44 0.92 ;
        RECT 1.36 0.52 1.54 0.73 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END OAI32X1

MACRO TLATNCAX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX6 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.35 3.32 1.38 ;
        RECT 3.26 0.6 3.34 0.81 ;
        RECT 3.67 0.35 3.73 1.38 ;
        RECT 3.26 0.75 4.14 0.81 ;
        RECT 4.08 0.35 4.14 1.38 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 0.92 0.68 1.085 ;
        RECT 0.6 1.005 0.765 1.085 ;
        RECT 0.685 1.005 0.765 1.335 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.775 0.5 0.895 ;
        RECT 0.42 0.725 0.5 1.04 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END TLATNCAX6

MACRO OA22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 1.39 1.54 1.49 ;
        RECT 1.46 1.36 1.655 1.42 ;
        RECT 1.595 0.425 1.655 1.42 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.76 1.14 1.26 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.56 0.73 ;
        RECT 0.48 0.6 0.56 1.08 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.98 0.74 1.11 ;
        RECT 0.72 0.67 0.8 1.06 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OA22XL

MACRO AND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X8 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.045 0.48 1.165 0.54 ;
        RECT 1.13 0.98 1.19 1.425 ;
        RECT 1.455 0.48 1.575 0.555 ;
        RECT 1.54 0.98 1.6 1.425 ;
        RECT 1.865 0.48 1.985 0.555 ;
        RECT 1.95 0.98 2.01 1.425 ;
        RECT 2.06 0.495 2.12 1.04 ;
        RECT 2.06 0.495 2.14 0.73 ;
        RECT 1.105 0.495 2.305 0.555 ;
        RECT 1.13 0.98 2.42 1.04 ;
        RECT 2.26 0.48 2.395 0.54 ;
        RECT 2.36 0.98 2.42 1.425 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.805 0.605 1.045 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.215 0.625 0.335 0.71 ;
        RECT 0.035 0.625 0.785 0.705 ;
        RECT 0.705 0.625 0.785 0.745 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END AND2X8

MACRO TLATNX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNX4 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.53 1.005 2.59 1.34 ;
        RECT 2.65 0.455 2.71 0.575 ;
        RECT 2.53 1.005 2.765 1.085 ;
        RECT 2.865 0.515 2.925 1.065 ;
        RECT 2.53 1.005 3 1.065 ;
        RECT 2.94 1.005 3 1.34 ;
        RECT 3.12 0.455 3.18 0.575 ;
        RECT 2.65 0.515 3.18 0.575 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.77 0.455 0.83 0.575 ;
        RECT 0.86 0.79 0.92 1.34 ;
        RECT 0.88 0.515 0.94 1.01 ;
        RECT 0.86 0.95 1.33 1.01 ;
        RECT 1.24 0.455 1.3 0.575 ;
        RECT 0.77 0.515 1.3 0.575 ;
        RECT 1.27 0.95 1.33 1.34 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.66 0.62 4.74 1.12 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.565 0.585 0.85 ;
        RECT 0.375 0.77 0.585 0.85 ;
        RECT 0.435 0.565 0.67 0.705 ;
    END
  END GN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.2 0.06 ;
    END
  END VSS
END TLATNX4

MACRO SMDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX8 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.86 0.695 6.92 0.945 ;
        RECT 6.8 0.885 6.92 0.945 ;
        RECT 6.86 0.695 7.08 0.755 ;
        RECT 7.035 0.625 7.205 0.705 ;
        RECT 7.02 0.645 7.715 0.705 ;
        RECT 7.655 0.645 7.715 0.765 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.18 0.805 7.375 1.01 ;
        RECT 7.18 0.805 7.555 0.885 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.46 0.535 6.54 0.995 ;
        RECT 6.42 0.885 6.54 0.995 ;
    END
  END D0
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.24 0.65 6.32 1.005 ;
        RECT 6.26 0.525 6.34 0.73 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.565 5.34 1.01 ;
        RECT 5.26 0.86 5.395 1.01 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.82 0.64 2.93 0.895 ;
        RECT 2.605 0.815 2.93 0.895 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.54 0.14 1.345 ;
        RECT 0.49 0.54 0.55 1.345 ;
        RECT 0.06 0.6 0.96 0.66 ;
        RECT 0.9 0.54 0.96 1.345 ;
        RECT 0.9 0.74 1.325 0.8 ;
        RECT 1.265 0.59 1.325 0.96 ;
        RECT 1.31 0.53 1.37 0.65 ;
        RECT 1.31 0.9 1.37 1.345 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8 0.06 ;
    END
  END VSS
END SMDFFHQX8

MACRO AOI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.56 0.36 0.62 0.48 ;
        RECT 0.56 0.42 0.94 0.48 ;
        RECT 0.88 0.42 0.94 1.44 ;
        RECT 0.88 0.6 1.14 0.73 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.56 0.34 1.06 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.58 0.56 1.06 ;
        RECT 0.46 0.79 0.56 1.06 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.58 0.74 1.04 ;
        RECT 0.66 0.58 0.78 0.66 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END AOI21X1

MACRO DFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRX4 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.07 0.485 5.14 1.29 ;
        RECT 5.06 0.79 5.14 1.29 ;
        RECT 5.06 0.9 5.55 0.96 ;
        RECT 5.49 0.9 5.55 1.29 ;
        RECT 5.07 0.485 5.66 0.545 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.79 4.32 1.29 ;
        RECT 4.28 0.485 4.34 0.96 ;
        RECT 4.26 0.9 4.73 0.96 ;
        RECT 4.13 0.485 4.72 0.545 ;
        RECT 4.67 0.9 4.73 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.125 0.625 1.42 0.895 ;
        RECT 1.125 0.815 1.435 0.895 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.69 0.405 1.055 ;
        RECT 0.325 0.79 0.54 1.055 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.98 0.14 1.11 ;
        RECT 0.095 0.695 0.225 1.055 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END DFFTRX4

MACRO TLATNCAX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX3 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.84 0.54 2.92 0.66 ;
        RECT 2.84 1.01 2.9 1.4 ;
        RECT 2.86 0.54 2.92 1.07 ;
        RECT 2.86 0.79 2.94 1.07 ;
        RECT 2.84 1.01 3.31 1.07 ;
        RECT 3.25 0.54 3.31 0.68 ;
        RECT 2.86 0.62 3.31 0.68 ;
        RECT 3.25 1.01 3.31 1.4 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.49 0.815 0.855 0.895 ;
        RECT 0.775 0.815 0.855 1.03 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.06 0.46 0.23 0.54 ;
        RECT 0.15 0.46 0.23 0.82 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END TLATNCAX3

MACRO FILL4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL4 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.8 0.06 ;
    END
  END VSS
END FILL4

MACRO OAI31XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.795 1.21 0.855 1.33 ;
        RECT 0.84 0.98 0.9 1.27 ;
        RECT 1.08 0.255 1.14 1.11 ;
        RECT 0.84 0.98 1.14 1.11 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 1.1 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.9 0.42 0.98 0.88 ;
        RECT 0.86 0.6 0.98 0.88 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.61 0.74 1.11 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END OAI31XL

MACRO NOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X1 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.49 0.52 0.63 ;
        RECT 0.46 0.57 0.72 0.63 ;
        RECT 0.66 0.57 0.72 1.29 ;
        RECT 0.66 0.6 0.74 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.57 0.34 1.07 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.98 0.54 1.21 ;
        RECT 0.48 0.73 0.56 1.085 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.8 0.06 ;
    END
  END VSS
END NOR2X1

MACRO SDFFSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX4 0 0 ;
  SIZE 9.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.275 0.915 8.335 1.305 ;
        RECT 8.275 0.915 8.38 0.975 ;
        RECT 8.32 0.45 8.385 0.92 ;
        RECT 8.32 0.79 8.54 0.92 ;
        RECT 8.32 0.86 8.7 0.92 ;
        RECT 8.64 0.86 8.7 1.015 ;
        RECT 8.685 0.955 8.745 1.305 ;
        RECT 8.265 0.45 8.855 0.51 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.415 0.915 7.475 1.305 ;
        RECT 7.48 0.45 7.54 0.975 ;
        RECT 7.46 0.79 7.54 0.975 ;
        RECT 7.415 0.915 7.885 0.975 ;
        RECT 7.825 0.915 7.885 1.305 ;
        RECT 7.325 0.45 7.915 0.51 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.575 0.555 4.655 0.895 ;
        RECT 4.575 0.815 4.815 0.895 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.31 0.555 4.39 0.895 ;
        RECT 4.235 0.815 4.475 0.895 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 0.625 1.535 0.895 ;
        RECT 1.455 0.625 1.765 0.705 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.185 0.585 1.265 0.805 ;
        RECT 1.26 0.725 1.34 1.01 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.2 0.805 0.365 0.98 ;
        RECT 0.2 0.9 0.605 0.98 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 0.585 0.36 0.705 ;
        RECT 0.62 0.26 0.68 0.705 ;
        RECT 0.3 0.585 0.68 0.645 ;
        RECT 0.62 0.625 0.765 0.705 ;
        RECT 0.62 0.26 1.085 0.32 ;
        RECT 1.025 0.26 1.085 0.965 ;
        RECT 1.025 0.905 1.145 0.965 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 9.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 9.6 0.06 ;
    END
  END VSS
END SDFFSRX4

MACRO SMDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX2 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.54 0.34 0.92 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.295 0.875 0.355 1.31 ;
    END
  END Q
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.46 0.695 5.52 0.945 ;
        RECT 5.4 0.885 5.52 0.945 ;
        RECT 5.46 0.695 5.735 0.755 ;
        RECT 5.675 0.645 6.315 0.705 ;
        RECT 6.035 0.625 6.315 0.705 ;
        RECT 6.255 0.625 6.315 0.745 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.835 0.805 6.155 1.01 ;
        RECT 5.78 0.885 6.155 1.01 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.545 5.14 0.93 ;
        RECT 4.945 0.85 5.14 0.93 ;
    END
  END D0
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.765 0.65 4.845 0.945 ;
        RECT 4.86 0.54 4.94 0.73 ;
        RECT 4.765 0.65 4.94 0.73 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.79 3.74 0.92 ;
        RECT 3.84 0.65 3.92 0.92 ;
        RECT 3.66 0.84 3.92 0.92 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.75 0.74 1.25 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.6 0.06 ;
    END
  END VSS
END SMDFFHQX2

MACRO MX4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.08 0.41 0.14 0.85 ;
        RECT 0.1 0.79 0.16 1.375 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.445 0.835 3.565 0.905 ;
        RECT 3.505 0.835 3.565 1.405 ;
        RECT 2.405 1.345 3.565 1.405 ;
        RECT 4.035 0.815 4.165 0.895 ;
        RECT 3.445 0.835 4.165 0.895 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.465 0.625 3.765 0.705 ;
        RECT 3.615 0.655 3.935 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.885 0.805 2.965 1.085 ;
        RECT 2.835 1.005 3.135 1.085 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.655 0.805 2.735 1.085 ;
        RECT 2.435 1.005 2.735 1.085 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.82 0.625 1.965 0.705 ;
        RECT 1.885 0.625 1.965 1.01 ;
        RECT 1.885 0.835 2.015 1.01 ;
    END
  END D
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 0.625 0.565 0.705 ;
        RECT 0.505 0.645 0.625 0.98 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END MX4X1

MACRO NOR3BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.43 0.14 1.27 ;
        RECT 0.13 0.37 0.19 0.51 ;
        RECT 0.08 1.21 0.305 1.27 ;
        RECT 0.245 1.21 0.305 1.33 ;
        RECT 0.54 0.37 0.6 0.51 ;
        RECT 0.08 0.45 0.6 0.51 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.645 0.94 1.145 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END NOR3BX1

MACRO SDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX1 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.54 0.92 1.315 ;
        RECT 0.86 0.6 0.94 0.73 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.28 0.73 ;
        RECT 0.2 0.54 0.28 1.29 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.38 0.64 4.44 0.965 ;
        RECT 4.32 0.905 4.44 0.965 ;
        RECT 4.38 0.64 5.165 0.7 ;
        RECT 4.93 0.585 4.99 0.705 ;
        RECT 4.93 0.625 5.165 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.835 0.805 5.21 0.935 ;
        RECT 4.76 0.855 5.21 0.935 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.585 3.94 0.73 ;
        RECT 3.86 0.65 4.06 0.73 ;
        RECT 3.98 0.65 4.06 0.965 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.19 0.88 1.27 1.085 ;
        RECT 1.035 1.005 1.27 1.085 ;
        RECT 1.2 0.75 1.28 0.96 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END SDFFX1

MACRO AND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X6 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.08 0.275 1.14 0.585 ;
        RECT 1.095 0.9 1.155 1.37 ;
        RECT 1.49 0.275 1.55 0.585 ;
        RECT 1.505 0.9 1.565 1.37 ;
        RECT 1.66 0.525 1.72 0.96 ;
        RECT 1.66 0.79 1.74 0.96 ;
        RECT 1.095 0.9 1.975 0.96 ;
        RECT 1.9 0.275 1.96 0.585 ;
        RECT 1.08 0.525 1.96 0.585 ;
        RECT 1.915 0.9 1.975 1.37 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 0.785 0.565 0.99 ;
        RECT 0.285 0.785 0.66 0.865 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.035 0.625 0.185 0.715 ;
        RECT 0.125 0.625 0.185 0.78 ;
        RECT 0.035 0.625 0.82 0.685 ;
        RECT 0.76 0.625 0.82 0.755 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END AND2X6

MACRO SEDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX8 0 0 ;
  SIZE 8.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.76 0.635 7.82 1.01 ;
        RECT 8.035 0.625 8.165 0.705 ;
        RECT 7.76 0.635 8.165 0.695 ;
        RECT 8.035 0.645 8.61 0.705 ;
        RECT 8.55 0.645 8.61 0.765 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.14 0.805 8.45 0.895 ;
        RECT 8.37 0.805 8.45 1.075 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.62 7.34 1.12 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.085 0.64 6.165 0.95 ;
        RECT 6.035 0.815 6.165 0.95 ;
        RECT 6.085 0.64 6.305 0.72 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.585 0.7 2.74 0.92 ;
        RECT 2.66 0.7 2.74 1.125 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.54 0.14 1.345 ;
        RECT 0.06 0.645 0.55 0.705 ;
        RECT 0.49 0.54 0.55 1.345 ;
        RECT 0.9 0.54 0.96 1.345 ;
        RECT 0.49 0.74 1.325 0.8 ;
        RECT 1.265 0.585 1.325 0.96 ;
        RECT 1.31 0.525 1.37 0.645 ;
        RECT 1.31 0.9 1.37 1.345 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.8 0.06 ;
    END
  END VSS
END SEDFFHQX8

MACRO DFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.6 4.17 0.73 ;
        RECT 4.09 0.57 4.17 0.94 ;
        RECT 4.11 0.88 4.19 1.29 ;
        RECT 4.09 0.57 4.25 0.65 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.57 3.78 0.73 ;
        RECT 3.72 0.57 3.78 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.535 3.34 0.895 ;
        RECT 3.18 0.77 3.4 0.895 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.575 0.2 0.73 ;
        RECT 0.12 0.575 0.2 1.015 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END DFFTRX2

MACRO TLATNTSCAX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX4 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.575 1.005 0.815 1.175 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.815 0.925 0.905 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.98 0.14 1.15 ;
        RECT 0.095 0.685 0.175 1.06 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.445 0.465 3.52 0.585 ;
        RECT 3.445 0.97 3.505 1.385 ;
        RECT 3.46 0.465 3.52 0.73 ;
        RECT 3.46 0.6 3.54 0.73 ;
        RECT 3.49 0.67 3.55 1.03 ;
        RECT 3.46 0.67 3.915 0.73 ;
        RECT 3.855 0.465 3.915 1.385 ;
    END
  END ECK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.2 0.06 ;
    END
  END VSS
END TLATNTSCAX4

MACRO DFFQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX4 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.485 0.675 3.565 0.975 ;
        RECT 3.485 0.815 3.765 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.46 0.34 0.96 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 0.485 0.72 0.545 ;
        RECT 0.66 0.485 0.72 1.355 ;
        RECT 0.66 0.6 0.74 0.73 ;
        RECT 0.66 0.67 1.105 0.73 ;
        RECT 1.045 0.485 1.105 1.02 ;
        RECT 1.07 0.965 1.13 1.355 ;
        RECT 1.045 0.485 1.185 0.545 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.2 0.06 ;
    END
  END VSS
END DFFQX4

MACRO AND3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X8 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.62 0.93 1.68 1.375 ;
        RECT 1.59 0.57 1.71 0.63 ;
        RECT 2.03 0.93 2.09 1.375 ;
        RECT 2 0.57 2.12 0.645 ;
        RECT 2.44 0.93 2.5 1.375 ;
        RECT 2.41 0.57 2.53 0.645 ;
        RECT 2.66 0.585 2.72 0.99 ;
        RECT 2.66 0.585 2.74 0.73 ;
        RECT 1.62 0.93 2.91 0.99 ;
        RECT 1.665 0.585 2.85 0.645 ;
        RECT 2.85 0.93 2.91 1.375 ;
        RECT 2.805 0.57 2.94 0.63 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.63 0.815 0.86 0.995 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.655 1.14 0.715 ;
        RECT 1.06 0.655 1.14 0.92 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.495 0.34 0.76 ;
        RECT 0.26 0.6 0.34 0.76 ;
        RECT 0.28 0.495 1.33 0.555 ;
        RECT 1.27 0.495 1.33 0.735 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END AND3X8

MACRO AOI221X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 0.4 0.92 0.46 ;
        RECT 1.46 0.22 1.54 0.48 ;
        RECT 0.87 0.42 1.54 0.48 ;
        RECT 1.48 0.22 1.54 1.46 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.58 0.94 1.08 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.58 1.14 1.08 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.45 0.34 0.95 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.58 1.34 1.04 ;
        RECT 1.26 0.65 1.38 0.73 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.54 0.72 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END AOI221X1

MACRO TLATNX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNX2 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.6 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.6 1.71 ;
    END
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.685 0.515 0.895 ;
        RECT 0.195 0.815 0.515 0.895 ;
        RECT 0.435 0.685 0.565 0.765 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.625 1.975 0.895 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.46 2.34 1.29 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.105 0.46 3.185 1.29 ;
        RECT 3.105 0.625 3.365 0.705 ;
    END
  END Q
END TLATNX2

MACRO INVXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVXL 0 0 ;
  SIZE 0.40 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 0.9 0.375 0.98 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.72 0.195 0.8 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.40 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.40 0.06 ;
    END
  END VSS
END INVXL

MACRO ADDFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFXL 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.295 3.92 1.2 ;
        RECT 3.86 0.6 3.94 0.73 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.48 0.14 0.92 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.06 0.86 0.375 0.92 ;
        RECT 0.315 0.285 0.375 0.54 ;
        RECT 0.08 0.48 0.375 0.54 ;
        RECT 0.315 0.86 0.375 1.045 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.055 0.785 1.115 0.905 ;
        RECT 1.58 0.845 1.765 1.085 ;
        RECT 1.055 0.845 2.03 0.905 ;
        RECT 1.97 0.82 3.36 0.88 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.83 0.67 0.955 0.73 ;
        RECT 0.895 0.625 1.235 0.685 ;
        RECT 1.185 0.66 3.54 0.705 ;
        RECT 0.895 0.645 1.395 0.685 ;
        RECT 1.335 0.66 3.54 0.72 ;
        RECT 3.46 0.66 3.54 1.005 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.495 0.435 1.765 0.56 ;
        RECT 1.495 0.5 3.15 0.56 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END ADDFXL

MACRO INVX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX6 0 0 ;
  SIZE 1.20 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.075 0.70 1.155 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.72 0.15 0.87 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.20 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.20 0.06 ;
    END
  END VSS
END INVX6

MACRO XNOR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3XL 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.24 0.57 4.365 0.705 ;
        RECT 4.235 0.625 4.365 0.705 ;
        RECT 4.305 0.57 4.365 1.1 ;
        RECT 4.24 1.04 4.365 1.1 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.175 0.92 ;
        RECT 0.095 0.635 0.175 1.1 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.625 0.515 0.78 ;
        RECT 0.46 0.7 0.54 1.1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.925 0.665 3.095 0.725 ;
        RECT 3.035 0.665 3.095 0.935 ;
        RECT 3.035 0.815 3.165 0.935 ;
        RECT 3.035 0.875 3.365 0.935 ;
    END
  END C
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END XNOR3XL

MACRO OR4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.4 1.74 1.355 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 0.73 ;
        RECT 0.66 0.6 0.92 0.68 ;
        RECT 0.84 0.48 0.92 0.75 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.48 0.56 0.96 ;
        RECT 0.46 0.79 0.56 0.96 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.48 0.36 0.96 ;
        RECT 0.26 0.79 0.36 0.96 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.195 0.35 1.275 0.76 ;
        RECT 1.195 0.625 1.365 0.705 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END OR4X2

MACRO AO21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.08 0.37 1.14 0.54 ;
        RECT 1.06 0.41 1.14 0.54 ;
        RECT 1.06 0.48 1.28 0.54 ;
        RECT 1.22 0.48 1.28 1.48 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.45 0.34 0.95 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.54 0.72 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.61 0.73 0.91 ;
        RECT 0.66 0.79 0.74 1.1 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END AO21X1

MACRO OAI221XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 1.115 0.985 1.3 ;
        RECT 1.645 0.325 1.705 1.3 ;
        RECT 0.925 1.115 1.705 1.175 ;
        RECT 1.56 1.17 1.74 1.3 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.675 0.34 1.175 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 0.815 1.145 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 1.17 0.54 1.3 ;
        RECT 0.465 0.805 0.545 1.25 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.515 1.34 1.015 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.52 1.545 1.015 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OAI221XL

MACRO NOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 0.35 0.51 0.63 ;
        RECT 0.45 0.57 0.92 0.63 ;
        RECT 0.86 0.49 0.92 1.29 ;
        RECT 0.86 0.79 0.94 0.92 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.98 0.74 1.21 ;
        RECT 0.68 0.73 0.76 1.11 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.57 0.34 1.07 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.73 0.54 1.23 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END NOR3X1

MACRO AND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X4 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 1.09 1.035 1.48 ;
        RECT 0.945 0.42 1.065 0.48 ;
        RECT 1.015 0.44 1.52 0.5 ;
        RECT 1.4 0.38 1.46 0.5 ;
        RECT 1.4 1.09 1.46 1.48 ;
        RECT 1.46 0.44 1.52 1.15 ;
        RECT 0.975 1.09 1.52 1.15 ;
        RECT 1.46 0.6 1.54 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.76 0.74 1.26 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.06 0.625 0.4 0.705 ;
        RECT 0.32 0.625 0.4 0.815 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END AND2X4

MACRO TLATNCAX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX12 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.61 0.26 0.67 0.57 ;
        RECT 0.61 0.9 0.67 1.02 ;
        RECT 0.99 0.51 1.05 0.99 ;
        RECT 1.02 0.26 1.08 0.57 ;
        RECT 0.99 0.79 1.14 0.99 ;
        RECT 0.61 0.9 1.14 0.99 ;
        RECT 1.43 0.26 1.49 0.57 ;
        RECT 1.84 0.26 1.9 0.57 ;
        RECT 2.25 0.26 2.31 0.57 ;
        RECT 0.61 0.51 2.31 0.57 ;
        RECT 0.61 0.93 2.34 0.99 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.13 0.85 5.21 1.06 ;
        RECT 5.13 0.98 5.34 1.06 ;
        RECT 5.26 0.98 5.34 1.22 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.62 0.325 0.7 ;
        RECT 0.235 0.62 0.325 0.895 ;
        RECT 0.235 0.815 0.51 0.895 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END TLATNCAX12

MACRO XOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.5 0.32 1.465 ;
        RECT 0.26 0.98 0.335 1.465 ;
        RECT 0.26 0.98 0.34 1.135 ;
        RECT 0.245 0.5 0.365 0.56 ;
        RECT 0.26 1.075 0.7 1.135 ;
        RECT 0.64 0.39 0.7 0.61 ;
        RECT 0.26 0.55 0.7 0.61 ;
        RECT 0.64 1.075 0.7 1.405 ;
        RECT 0.685 0.33 0.745 0.45 ;
        RECT 0.685 1.345 0.745 1.465 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.745 0.625 2.205 0.705 ;
        RECT 2.125 0.625 2.205 0.745 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.96 0.71 1.165 1.085 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END XOR2X4

MACRO SDFFSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX1 0 0 ;
  SIZE 7 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.98 1.14 1.11 ;
        RECT 1.08 0.9 1.14 1.29 ;
        RECT 1.08 0.9 1.255 1.04 ;
        RECT 1.195 0.54 1.255 1.04 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.57 0.54 0.65 ;
        RECT 0.42 0.9 0.5 1.29 ;
        RECT 0.46 0.57 0.54 0.98 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.075 0.655 6.135 0.93 ;
        RECT 6.015 0.87 6.135 0.93 ;
        RECT 6.355 0.585 6.415 0.715 ;
        RECT 6.075 0.655 6.495 0.715 ;
        RECT 6.355 0.625 6.565 0.705 ;
        RECT 6.355 0.645 6.725 0.705 ;
        RECT 6.665 0.585 6.725 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.235 0.815 6.695 0.895 ;
        RECT 6.46 0.815 6.695 0.935 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.46 0.515 5.54 0.8 ;
        RECT 5.46 0.72 5.755 0.8 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.55 5.36 0.73 ;
        RECT 5.28 0.515 5.36 0.995 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.325 2.295 0.895 ;
        RECT 2.235 0.815 2.365 0.895 ;
        RECT 1.855 0.835 2.365 0.895 ;
        RECT 2.235 0.325 3.075 0.385 ;
        RECT 3.015 0.35 3.455 0.41 ;
        RECT 3.395 0.33 3.515 0.39 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7 0.06 ;
    END
  END VSS
END SDFFSX1

MACRO AOI2BB2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X4 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.4 0.445 1.52 0.505 ;
        RECT 2.02 0.445 2.14 0.525 ;
        RECT 2.475 0.465 2.535 0.865 ;
        RECT 2.475 0.805 2.695 0.865 ;
        RECT 2.635 0.805 2.695 1.085 ;
        RECT 1.47 0.465 2.7 0.525 ;
        RECT 2.665 0.995 2.765 1.115 ;
        RECT 2.65 0.445 2.99 0.505 ;
        RECT 3.075 0.995 3.135 1.115 ;
        RECT 3.485 0.995 3.545 1.115 ;
        RECT 3.66 0.445 3.785 0.505 ;
        RECT 3.725 0.445 3.785 1.055 ;
        RECT 2.635 0.995 3.955 1.055 ;
        RECT 3.895 0.995 3.955 1.115 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 0.815 3.625 0.895 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.635 0.625 2.765 0.705 ;
        RECT 3.5 0.285 3.56 0.705 ;
        RECT 2.635 0.645 3.56 0.705 ;
        RECT 3.5 0.285 3.945 0.345 ;
        RECT 3.885 0.285 3.945 0.7 ;
        RECT 3.885 0.64 4.06 0.7 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.695 0.54 1.195 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.695 0.34 1.195 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END AOI2BB2X4

MACRO NOR4BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.45 0.14 1.27 ;
        RECT 0.08 1.21 0.5 1.27 ;
        RECT 0.44 1.21 0.5 1.425 ;
        RECT 0.545 0.37 0.605 0.51 ;
        RECT 0.92 0.4 1.03 0.46 ;
        RECT 0.08 0.45 0.98 0.51 ;
        RECT 0.97 0.34 1.03 0.46 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.61 1.54 1.11 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.865 0.81 1.36 0.89 ;
        RECT 1.035 0.81 1.36 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.635 0.765 1.085 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END NOR4BX1

MACRO SEDFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX1 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.42 0.54 5.5 1.08 ;
        RECT 5.315 1 5.5 1.08 ;
        RECT 5.42 0.6 5.54 0.73 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.54 0.14 1.29 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.86 0.98 7.94 1.17 ;
        RECT 7.89 0.7 7.97 1.06 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.985 0.77 7.54 0.85 ;
        RECT 7.46 0.77 7.54 0.92 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.86 0.875 5.94 1.205 ;
        RECT 5.86 0.875 6.11 0.955 ;
    END
  END RN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.08 0.64 4.16 0.96 ;
        RECT 4.08 0.64 4.34 0.92 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.835 0.625 3.98 0.705 ;
        RECT 3.92 0.48 3.98 0.82 ;
        RECT 3.92 0.48 4.66 0.54 ;
        RECT 4.6 0.48 4.66 0.82 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.67 3.35 1.12 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.2 0.06 ;
    END
  END VSS
END SEDFFTRX1

MACRO SEDFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX4 0 0 ;
  SIZE 9.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.905 0.49 5.965 1.085 ;
        RECT 5.705 1.025 5.965 1.085 ;
        RECT 5.835 1.005 6.17 1.065 ;
        RECT 6.11 1.025 6.295 1.085 ;
        RECT 5.835 0.49 6.425 0.55 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.46 5.12 1.085 ;
        RECT 4.735 1.025 5.165 1.085 ;
        RECT 5.035 1.005 5.325 1.065 ;
        RECT 5.265 1.005 5.325 1.125 ;
        RECT 4.895 0.46 5.485 0.52 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9.26 0.41 9.34 0.91 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.86 0.79 8.95 0.92 ;
        RECT 8.87 0.74 8.95 0.92 ;
        RECT 8.43 0.84 8.95 0.92 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.78 7.39 1.23 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.4 0.65 4.54 0.73 ;
        RECT 4.46 0.6 4.54 1.04 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.19 0.805 0.58 0.985 ;
        RECT 0.19 0.905 0.59 0.985 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.225 0.625 0.365 0.705 ;
        RECT 0.545 0.3 0.605 0.705 ;
        RECT 0.225 0.645 0.75 0.705 ;
        RECT 0.545 0.3 1.07 0.36 ;
        RECT 1.01 0.3 1.07 0.85 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 9.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 9.6 0.06 ;
    END
  END VSS
END SEDFFTRX4

MACRO NAND3BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.44 0.14 1.26 ;
        RECT 0.06 0.98 0.14 1.26 ;
        RECT 0.145 1.2 0.205 1.48 ;
        RECT 0.2 0.38 0.26 0.5 ;
        RECT 0.08 0.44 0.26 0.5 ;
        RECT 0.06 1.2 0.615 1.26 ;
        RECT 0.555 1.2 0.615 1.48 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.76 0.94 1.26 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.54 1.1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END NAND3BX1

MACRO DFFQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX2 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.79 3.12 1.355 ;
        RECT 3.08 0.54 3.14 0.92 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.59 0.94 0.73 ;
        RECT 0.86 0.65 1.055 0.73 ;
        RECT 0.975 0.65 1.055 0.975 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.06 0.625 0.37 0.73 ;
        RECT 0.29 0.625 0.37 0.87 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END DFFQX2

MACRO AND3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X6 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 0.345 1.66 0.655 ;
        RECT 1.6 0.92 1.66 1.37 ;
        RECT 2.01 0.345 2.07 0.655 ;
        RECT 2.01 0.92 2.07 1.37 ;
        RECT 2.26 0.595 2.32 0.98 ;
        RECT 2.26 0.79 2.34 0.98 ;
        RECT 1.6 0.92 2.48 0.98 ;
        RECT 2.42 0.345 2.48 0.655 ;
        RECT 1.6 0.595 2.48 0.655 ;
        RECT 2.42 0.92 2.48 1.37 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.53 0.815 0.96 0.965 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.47 0.655 1.14 0.715 ;
        RECT 1.06 0.655 1.14 0.92 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.37 0.73 ;
        RECT 0.31 0.495 0.37 0.735 ;
        RECT 0.31 0.495 1.32 0.555 ;
        RECT 1.26 0.495 1.32 0.75 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.6 0.06 ;
    END
  END VSS
END AND3X6

MACRO AOI221X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.76 0.445 0.88 0.505 ;
        RECT 1.38 0.445 1.5 0.525 ;
        RECT 1.835 0.625 1.965 0.705 ;
        RECT 1.905 0.465 1.965 1.055 ;
        RECT 2.37 0.445 2.49 0.525 ;
        RECT 3.135 0.445 3.255 0.525 ;
        RECT 3.675 0.445 3.795 0.525 ;
        RECT 3.835 0.995 3.895 1.135 ;
        RECT 0.83 0.465 4.165 0.525 ;
        RECT 4.115 0.445 4.235 0.505 ;
        RECT 1.905 0.995 4.305 1.055 ;
        RECT 4.245 0.995 4.305 1.135 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.815 1.425 0.895 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.5 0.815 3.18 0.895 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.365 0.705 ;
        RECT 0.23 0.645 1.735 0.705 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.425 0.655 3.485 0.895 ;
        RECT 2.09 0.655 3.545 0.715 ;
        RECT 3.425 0.815 3.565 0.895 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.835 0.625 3.965 0.895 ;
        RECT 3.835 0.63 4.195 0.71 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END AOI221X4

MACRO XOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.28 0.495 0.34 1.215 ;
        RECT 0.28 1.155 0.435 1.215 ;
        RECT 0.375 0.435 0.435 0.555 ;
        RECT 0.28 0.495 0.435 0.555 ;
        RECT 0.375 1.155 0.435 1.275 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.825 1.565 0.885 ;
        RECT 1.435 0.815 1.565 0.895 ;
        RECT 1.335 0.815 1.785 0.875 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 0.815 0.8 0.895 ;
        RECT 0.72 0.815 0.8 1.195 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END XOR2X2

MACRO DFFRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX4 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.055 1.05 5.115 1.33 ;
        RECT 5.065 0.57 5.14 1.11 ;
        RECT 5.06 0.98 5.14 1.11 ;
        RECT 5.43 1.065 5.525 1.13 ;
        RECT 5.055 1.05 5.49 1.11 ;
        RECT 5.465 1.065 5.525 1.33 ;
        RECT 5.065 0.57 5.655 0.63 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.215 0.94 4.275 1.33 ;
        RECT 4.26 0.55 4.32 1 ;
        RECT 4.26 0.79 4.34 1 ;
        RECT 4.215 0.94 4.685 1 ;
        RECT 4.625 0.94 4.685 1.33 ;
        RECT 4.125 0.55 4.715 0.61 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.625 2.4 0.705 ;
        RECT 2.34 0.3 2.4 0.87 ;
        RECT 1.845 0.81 2.4 0.87 ;
        RECT 2.34 0.3 3.08 0.36 ;
        RECT 3.02 0.3 3.08 0.47 ;
        RECT 3.02 0.41 3.37 0.47 ;
        RECT 3.31 0.41 3.37 0.63 ;
        RECT 3.31 0.57 3.905 0.63 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.785 0.94 1.2 ;
        RECT 0.86 0.785 1.025 0.865 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.17 0.53 0.25 0.87 ;
        RECT 0.06 0.79 0.25 0.87 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END DFFRX4

MACRO AND4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X8 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.065 0.48 2.2 0.54 ;
        RECT 2.215 0.9 2.275 1.345 ;
        RECT 2.475 0.48 2.595 0.555 ;
        RECT 2.625 0.9 2.685 1.345 ;
        RECT 2.885 0.48 3.005 0.555 ;
        RECT 3.035 0.9 3.095 1.345 ;
        RECT 3.06 0.495 3.12 0.96 ;
        RECT 3.06 0.79 3.14 0.96 ;
        RECT 2.14 0.495 3.34 0.555 ;
        RECT 3.28 0.48 3.415 0.54 ;
        RECT 2.215 0.9 3.505 0.96 ;
        RECT 3.445 0.9 3.505 1.345 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.82 0.32 1.185 ;
        RECT 1.66 0.98 1.805 1.185 ;
        RECT 1.745 0.82 1.805 1.185 ;
        RECT 0.26 1.125 1.805 1.185 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 0.835 0.54 0.895 ;
        RECT 0.46 0.79 0.54 1.025 ;
        RECT 1.5 0.76 1.56 1.025 ;
        RECT 0.46 0.965 1.56 1.025 ;
        RECT 1.5 0.76 1.645 0.88 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.625 1.38 0.705 ;
        RECT 1.32 0.625 1.38 0.865 ;
        RECT 0.67 0.805 1.38 0.865 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.4 0.94 0.705 ;
        RECT 0.86 0.625 1.135 0.705 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.6 0.06 ;
    END
  END VSS
END AND4X8

MACRO SDFFRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRXL 0 0 ;
  SIZE 6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.47 0.92 1.385 ;
        RECT 0.86 0.98 0.94 1.385 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.285 0.73 ;
        RECT 0.205 0.54 0.285 1.02 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.805 0.465 4.865 0.91 ;
        RECT 5.07 0.465 5.13 0.725 ;
        RECT 4.805 0.465 5.695 0.525 ;
        RECT 5.635 0.465 5.695 0.705 ;
        RECT 5.635 0.625 5.765 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.23 0.625 5.365 0.9 ;
        RECT 5.23 0.82 5.535 0.9 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.79 4.54 0.99 ;
        RECT 4.465 0.495 4.545 0.87 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.815 1.765 0.92 ;
        RECT 1.635 0.82 2.11 0.9 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.98 1.14 1.26 ;
        RECT 1.13 0.83 1.21 1.085 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6 0.06 ;
    END
  END VSS
END SDFFRXL

MACRO SDFFNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX1 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.89 0.555 0.95 1.11 ;
        RECT 0.86 0.98 0.95 1.11 ;
        RECT 0.935 1.035 0.995 1.425 ;
        RECT 0.94 0.515 1 0.635 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.29 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.235 0.625 7.365 0.725 ;
        RECT 7.04 0.645 7.52 0.725 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.2 0.825 7.52 1.085 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.48 0.67 6.56 1.15 ;
        RECT 6.46 0.98 6.56 1.15 ;
    END
  END D
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.67 6.36 0.92 ;
        RECT 6.28 0.67 6.36 1.15 ;
    END
  END CKN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.815 2.365 0.895 ;
        RECT 2.13 0.835 2.365 0.895 ;
        RECT 2.305 0.815 2.365 0.985 ;
        RECT 2.305 0.925 3.22 0.985 ;
        RECT 3.16 0.925 3.22 1.235 ;
        RECT 3.16 1.175 4.12 1.235 ;
        RECT 4.06 1.175 4.12 1.405 ;
        RECT 4.06 1.345 4.515 1.405 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 0.895 1.365 1.205 ;
        RECT 1.095 1.005 1.365 1.205 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.8 0.06 ;
    END
  END VSS
END SDFFNSRX1

MACRO AOI31X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.73 0.37 0.79 0.51 ;
        RECT 0.73 0.45 1.12 0.51 ;
        RECT 1.06 0.45 1.12 1.48 ;
        RECT 1.06 0.6 1.14 0.73 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.45 0.34 0.95 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.61 0.94 1.11 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.61 0.73 1.1 ;
        RECT 0.65 0.61 0.74 0.92 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.54 0.35 ;
        RECT 0.47 0.27 0.55 0.71 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END AOI31X1

MACRO SDFFNSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX4 0 0 ;
  SIZE 9.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.045 0.915 8.105 1.305 ;
        RECT 8.08 0.48 8.14 0.975 ;
        RECT 8.06 0.79 8.14 0.975 ;
        RECT 8.045 0.915 8.515 0.975 ;
        RECT 8.455 0.915 8.515 1.305 ;
        RECT 8.08 0.48 8.67 0.54 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.48 7.32 1.305 ;
        RECT 7.225 0.915 7.32 1.305 ;
        RECT 7.26 0.79 7.34 0.92 ;
        RECT 7.26 0.86 7.695 0.92 ;
        RECT 7.635 0.86 7.695 1.305 ;
        RECT 7.14 0.48 7.73 0.54 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.035 0.625 4.165 0.705 ;
        RECT 4.085 0.655 4.59 0.735 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.635 0.625 3.935 0.705 ;
        RECT 3.855 0.625 3.935 0.905 ;
    END
  END SN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.7 1.54 1.2 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.65 1.34 1.15 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.715 0.54 1.075 ;
        RECT 0.46 0.715 0.68 0.92 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 0.555 0.36 0.675 ;
        RECT 0.66 0.41 0.84 0.615 ;
        RECT 0.3 0.555 0.84 0.615 ;
        RECT 0.78 0.295 0.84 0.795 ;
        RECT 0.78 0.295 1.16 0.355 ;
        RECT 1.1 0.295 1.16 1.06 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 9.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 9.4 0.06 ;
    END
  END VSS
END SDFFNSRX4

MACRO AND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X2 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.445 0.92 1.34 ;
        RECT 0.86 0.6 0.94 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.685 0.59 0.92 ;
        RECT 0.51 0.685 0.59 1.135 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.955 0.14 1.125 ;
        RECT 0.12 0.685 0.2 1.11 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END AND2X2

MACRO OR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.88 1.03 0.96 1.21 ;
        RECT 1.06 0.26 1.14 1.11 ;
        RECT 0.88 1.03 1.14 1.11 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 0.645 0.705 1.085 ;
        RECT 0.625 1.005 0.765 1.085 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.64 0.365 0.92 ;
        RECT 0.285 0.64 0.365 1.115 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.615 0.14 1.115 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OR3XL

MACRO CLKBUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX4 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.42 0.29 1.04 ;
        RECT 0.275 0.36 0.335 0.48 ;
        RECT 0.26 0.98 0.335 1.37 ;
        RECT 0.26 0.98 0.34 1.11 ;
        RECT 0.23 0.98 0.76 1.04 ;
        RECT 0.23 0.42 0.72 0.48 ;
        RECT 0.7 0.98 0.76 1.37 ;
        RECT 0.67 0.4 0.79 0.46 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.78 0.94 1.15 ;
        RECT 0.95 0.74 1.03 0.86 ;
        RECT 0.86 0.78 1.03 0.86 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END CLKBUFX4

MACRO AO22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 0.415 1.52 0.535 ;
        RECT 1.46 0.415 1.52 1.11 ;
        RECT 1.46 0.98 1.54 1.11 ;
        RECT 1.54 1.05 1.6 1.44 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 0.655 1.105 1.12 ;
        RECT 1.025 0.79 1.14 1 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.98 0.14 1.11 ;
        RECT 0.08 0.63 0.16 1.06 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.625 0.715 1.075 ;
        RECT 0.635 0.625 0.765 0.745 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.26 0.79 0.535 0.87 ;
        RECT 0.455 0.79 0.535 1.045 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END AO22X1

MACRO NOR4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 0.49 0.63 0.63 ;
        RECT 0.99 0.49 1.05 0.63 ;
        RECT 0.57 0.57 1.34 0.63 ;
        RECT 1.24 0.57 1.3 1.29 ;
        RECT 1.24 0.57 1.34 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.06 0.6 0.47 0.68 ;
        RECT 0.39 0.6 0.47 0.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.98 0.74 1.21 ;
        RECT 0.68 0.73 0.76 1.06 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.73 0.94 1.23 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.73 1.14 1.23 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END NOR4X1

MACRO NAND3BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX4 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.08 0.41 0.14 1.095 ;
        RECT 0.08 1.035 0.36 1.095 ;
        RECT 0.3 1.035 0.36 1.425 ;
        RECT 0.71 1.125 0.77 1.425 ;
        RECT 1.12 1.125 1.18 1.425 ;
        RECT 1.53 1.125 1.59 1.425 ;
        RECT 0.06 0.41 1.95 0.47 ;
        RECT 1.94 1.125 2 1.425 ;
        RECT 0.3 1.125 2.41 1.185 ;
        RECT 2.35 1.125 2.41 1.425 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.625 0.565 0.715 ;
        RECT 0.4 0.655 0.72 0.715 ;
        RECT 0.66 0.655 0.72 0.865 ;
        RECT 0.66 0.805 1.285 0.865 ;
        RECT 1.225 0.745 1.665 0.805 ;
        RECT 1.605 0.805 2.265 0.865 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.365 0.625 2.565 0.705 ;
        RECT 2.485 0.625 2.565 0.795 ;
        RECT 2.485 0.715 2.775 0.795 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 0.625 0.965 0.705 ;
        RECT 0.82 0.645 1.125 0.705 ;
        RECT 1.065 0.585 1.825 0.645 ;
        RECT 1.765 0.645 1.885 0.705 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3 0.06 ;
    END
  END VSS
END NAND3BX4

MACRO AND3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X4 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.895 0.57 1.015 0.63 ;
        RECT 1.04 1.08 1.1 1.47 ;
        RECT 1.335 0.57 1.525 0.65 ;
        RECT 0.965 0.59 1.525 0.65 ;
        RECT 1.45 1.08 1.51 1.47 ;
        RECT 1.465 0.57 1.525 1.14 ;
        RECT 1.04 1.08 1.525 1.14 ;
        RECT 1.465 0.79 1.74 0.92 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.91 0.78 1.06 ;
        RECT 0.7 0.98 0.94 1.06 ;
        RECT 0.86 0.98 0.94 1.25 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.26 0.65 0.44 0.73 ;
        RECT 0.36 0.65 0.44 1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.59 0.14 1.09 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END AND3X4

MACRO DFFRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX1 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.435 0.14 0.995 ;
        RECT 0.06 0.915 0.225 0.995 ;
        RECT 0.09 0.385 0.17 0.505 ;
        RECT 0.145 0.915 0.225 1.305 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.815 1.765 1.01 ;
        RECT 1.38 0.92 1.765 1.01 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.485 0.745 0.565 1.085 ;
        RECT 0.4 1.005 0.565 1.085 ;
        RECT 0.485 0.745 0.64 0.825 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.235 0.625 4.41 0.89 ;
        RECT 4.095 0.755 4.41 0.89 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END DFFRHQX1

MACRO AOI211XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 0.285 0.655 0.51 ;
        RECT 1.005 0.285 1.14 0.51 ;
        RECT 0.595 0.45 1.14 0.51 ;
        RECT 1.08 0.285 1.14 1.295 ;
        RECT 1.06 0.98 1.14 1.295 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.51 0.16 0.73 ;
        RECT 0.08 0.51 0.16 0.99 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 0.99 ;
        RECT 0.26 0.61 0.46 0.705 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.61 0.74 0.99 ;
        RECT 0.56 0.61 0.76 0.69 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.61 0.94 1.11 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END AOI211XL

MACRO DFFRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX2 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.31 0.565 4.37 0.975 ;
        RECT 4.36 0.915 4.42 1.305 ;
        RECT 4.31 0.565 4.45 0.625 ;
        RECT 4.36 0.915 4.54 1.11 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.535 3.92 1.305 ;
        RECT 3.86 0.925 3.94 1.11 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.455 0.89 3.535 1.085 ;
        RECT 3.375 1.005 3.76 1.085 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.815 1.365 0.895 ;
        RECT 1.285 0.855 1.695 0.935 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.365 0.815 0.445 1.185 ;
        RECT 0.235 1.005 0.445 1.185 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END DFFRX2

MACRO AND4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X6 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.245 0.275 2.305 0.585 ;
        RECT 2.45 0.9 2.51 1.37 ;
        RECT 2.655 0.275 2.715 0.585 ;
        RECT 2.86 0.525 2.92 1.37 ;
        RECT 2.86 0.79 2.94 1.37 ;
        RECT 3.065 0.275 3.125 0.585 ;
        RECT 2.245 0.525 3.125 0.585 ;
        RECT 2.45 0.9 3.33 0.96 ;
        RECT 3.27 0.9 3.33 1.37 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.395 0.82 0.455 1.185 ;
        RECT 1.86 0.82 1.92 1.185 ;
        RECT 0.395 1.125 1.92 1.185 ;
        RECT 1.86 0.82 1.94 1.11 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.835 0.74 0.895 ;
        RECT 0.66 0.79 0.74 1.025 ;
        RECT 1.7 0.845 1.76 1.025 ;
        RECT 0.66 0.965 1.76 1.025 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 0.625 1.515 0.865 ;
        RECT 0.84 0.805 1.515 0.865 ;
        RECT 1.435 0.625 1.565 0.705 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.41 0.94 0.685 ;
        RECT 0.86 0.605 1.165 0.685 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END AND4X6

MACRO OR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X4 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 0.855 1.035 1.405 ;
        RECT 0.945 0.4 1.065 0.46 ;
        RECT 1.015 0.42 1.52 0.48 ;
        RECT 0.975 0.855 1.52 0.915 ;
        RECT 1.4 0.36 1.46 0.48 ;
        RECT 1.4 1.015 1.46 1.405 ;
        RECT 1.46 0.42 1.52 1.075 ;
        RECT 1.46 0.6 1.54 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.605 0.74 0.74 0.86 ;
        RECT 0.66 0.74 0.74 1.185 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.06 0.6 0.345 0.68 ;
        RECT 0.265 0.6 0.345 0.845 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OR2X4

MACRO NAND4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.37 1.02 0.43 1.3 ;
        RECT 0.79 1.02 0.85 1.3 ;
        RECT 1.04 0.54 1.1 1.08 ;
        RECT 1.04 0.79 1.14 1.08 ;
        RECT 0.37 1.02 1.14 1.08 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.65 0.34 0.92 ;
        RECT 0.03 0.84 0.34 0.92 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.48 0.46 0.56 0.89 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.22 0.74 0.83 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.41 0.94 0.91 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END NAND4X1

MACRO AOI2BB2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X1 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 0.6 1.88 0.92 ;
        RECT 1.86 0.48 1.94 0.73 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.45 1.54 0.95 ;
    END
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.94 0.34 1.11 ;
        RECT 0.47 0.83 0.56 1.02 ;
        RECT 0.26 0.94 0.56 1.02 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.65 0.34 0.84 ;
        RECT 0.46 0.54 0.54 0.73 ;
        RECT 0.26 0.65 0.54 0.73 ;
    END
  END A1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.22 1.54 0.35 ;
        RECT 1.405 0.245 1.54 0.35 ;
        RECT 1.405 0.29 1.7 0.35 ;
        RECT 1.64 0.29 1.7 1.06 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END AOI2BB2X1

MACRO NAND2BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BXL 0 0 ;
  SIZE 1.00 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.04 0.72 0.135 0.8 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.72 0.9 0.8 1.095 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.865 0.31 0.945 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.00 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.00 0.06 ;
    END
  END VSS
END NAND2BXL

MACRO DFFSX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX4 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.54 5.32 1.33 ;
        RECT 5.26 0.6 5.34 1 ;
        RECT 5.26 0.94 5.73 1 ;
        RECT 5.67 0.94 5.73 1.33 ;
        RECT 5.73 0.54 5.79 0.66 ;
        RECT 5.26 0.6 5.79 0.66 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.32 0.505 4.38 0.625 ;
        RECT 4.44 0.94 4.5 1.33 ;
        RECT 4.46 0.565 4.52 1 ;
        RECT 4.46 0.79 4.54 1 ;
        RECT 4.44 0.94 4.91 1 ;
        RECT 4.79 0.505 4.85 0.625 ;
        RECT 4.32 0.565 4.85 0.625 ;
        RECT 4.85 0.94 4.91 1.33 ;
    END
  END Q
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.82 0.375 2 0.435 ;
        RECT 1.94 0.38 2.32 0.44 ;
        RECT 2.26 0.335 3.14 0.395 ;
        RECT 3.08 0.335 3.14 0.92 ;
        RECT 3.06 0.79 3.14 0.92 ;
        RECT 3.06 0.85 3.575 0.91 ;
        RECT 3.515 0.85 3.575 0.97 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.775 0.54 0.995 ;
        RECT 0.575 0.61 0.655 0.895 ;
        RECT 0.46 0.775 0.655 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.36 0.96 ;
        RECT 0.28 0.61 0.36 1.09 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END DFFSX4

MACRO OR3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X6 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.665 0.915 1.725 1.37 ;
        RECT 1.765 0.35 1.825 0.655 ;
        RECT 2.075 0.915 2.135 1.37 ;
        RECT 1.765 0.595 2.34 0.655 ;
        RECT 2.235 0.35 2.295 0.655 ;
        RECT 2.26 0.595 2.32 0.975 ;
        RECT 2.26 0.595 2.34 0.73 ;
        RECT 1.665 0.915 2.545 0.975 ;
        RECT 2.485 0.915 2.545 1.37 ;
        RECT 2.645 0.35 2.705 0.66 ;
        RECT 2.26 0.6 2.705 0.66 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.85 0.74 1.13 ;
        RECT 0.66 0.85 0.96 0.93 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.56 0.69 1.225 0.75 ;
        RECT 1.06 0.69 1.14 0.92 ;
        RECT 1.06 0.69 1.225 0.81 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.53 0.34 0.73 ;
        RECT 0.26 0.53 1.39 0.59 ;
        RECT 1.33 0.53 1.39 0.74 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END OR3X6

MACRO AND3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.145 0.48 1.205 0.66 ;
        RECT 1.145 0.6 1.34 0.66 ;
        RECT 1.26 0.6 1.32 1.42 ;
        RECT 1.26 0.6 1.34 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 1.005 0.915 1.455 ;
        RECT 0.835 1.005 0.965 1.085 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.56 0.34 0.73 ;
        RECT 0.26 0.56 0.575 0.64 ;
        RECT 0.495 0.56 0.575 0.735 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.56 0.16 1.04 ;
        RECT 0.06 0.79 0.16 1.04 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END AND3X2

MACRO ADDHXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHXL 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.465 2.72 0.585 ;
        RECT 2.66 0.98 2.74 1.135 ;
        RECT 2.71 0.525 2.77 1.04 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.435 0.34 1.23 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.79 0.74 1.135 ;
        RECT 0.785 0.76 0.865 0.91 ;
        RECT 0.66 0.79 0.865 0.91 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.56 0.73 ;
        RECT 0.66 0.305 0.72 0.66 ;
        RECT 0.46 0.6 0.72 0.66 ;
        RECT 0.66 0.305 1.345 0.365 ;
        RECT 1.285 0.305 1.345 0.72 ;
        RECT 1.605 0.305 1.665 0.72 ;
        RECT 1.285 0.66 1.665 0.72 ;
        RECT 1.605 0.305 1.725 0.365 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END ADDHXL

MACRO DFFRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.41 1.54 0.54 ;
        RECT 1.48 0.305 1.54 0.725 ;
        RECT 1.465 0.41 1.54 0.725 ;
        RECT 1.48 0.305 2 0.365 ;
        RECT 1.94 0.305 2 0.555 ;
        RECT 2.035 0.495 2.095 0.715 ;
        RECT 2.355 0.305 2.415 0.555 ;
        RECT 1.94 0.495 2.415 0.555 ;
        RECT 2.355 0.305 3.36 0.365 ;
        RECT 3.3 0.305 3.36 0.85 ;
        RECT 3.68 0.73 3.74 0.85 ;
        RECT 3.3 0.79 3.74 0.85 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.19 0.685 0.56 0.765 ;
        RECT 0.235 0.685 0.56 0.895 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.57 5.14 0.885 ;
        RECT 5.06 0.625 5.325 0.885 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.49 0.72 1.055 ;
        RECT 0.6 0.995 0.72 1.055 ;
        RECT 0.66 0.79 0.74 1.005 ;
        RECT 0.66 0.945 1.19 1.005 ;
        RECT 1.095 0.49 1.19 1.005 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END DFFRHQX4

MACRO NAND3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 1.105 0.94 1.165 ;
        RECT 0.87 0.54 0.94 1.225 ;
        RECT 0.86 0.98 0.94 1.225 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.395 0.74 0.88 ;
        RECT 0.66 0.76 0.755 0.88 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.03 0.735 0.11 1.005 ;
        RECT 0.03 0.79 0.34 1.005 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.48 0.48 0.56 0.89 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END NAND3XL

MACRO SEDFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFX4 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.205 0.485 6.265 0.625 ;
        RECT 6.26 0.565 6.32 1.11 ;
        RECT 6.26 0.98 6.34 1.11 ;
        RECT 6.045 1.05 6.34 1.11 ;
        RECT 6.26 1.005 6.575 1.065 ;
        RECT 6.515 1.02 6.635 1.08 ;
        RECT 6.615 0.485 6.675 0.625 ;
        RECT 6.205 0.565 6.675 0.625 ;
    END
  END QN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.045 0.795 7.105 0.955 ;
        RECT 7.29 0.725 7.35 0.855 ;
        RECT 7.045 0.795 7.35 0.855 ;
        RECT 7.46 0.6 7.54 0.785 ;
        RECT 7.29 0.725 7.74 0.785 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.44 0.98 7.54 1.11 ;
        RECT 7.45 0.885 7.795 1.085 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.83 0.725 5.91 1.195 ;
        RECT 5.83 0.725 5.94 0.925 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.635 0.51 4.765 0.59 ;
        RECT 4.685 0.51 4.765 0.96 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.435 0.69 4.575 0.98 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.54 0.335 1.345 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.26 0.67 0.7 0.73 ;
        RECT 0.64 0.6 0.7 0.975 ;
        RECT 0.685 0.54 0.745 0.66 ;
        RECT 0.685 0.915 0.745 1.345 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8 0.06 ;
    END
  END VSS
END SEDFFX4

MACRO AND4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 0.48 1.295 0.54 ;
        RECT 1.29 1.09 1.35 1.48 ;
        RECT 1.29 1.09 1.805 1.15 ;
        RECT 1.615 0.48 1.805 0.56 ;
        RECT 1.245 0.5 1.805 0.56 ;
        RECT 1.745 0.48 1.805 1.48 ;
        RECT 1.7 1.09 1.805 1.48 ;
        RECT 1.745 0.6 1.94 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.82 1.08 1.06 ;
        RECT 1.06 0.98 1.14 1.26 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.5 0.74 1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.52 0.56 0.74 ;
        RECT 0.48 0.52 0.56 1 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.99 ;
        RECT 0.28 0.51 0.36 0.73 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END AND4X4

MACRO OR4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X8 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.025 0.815 2.085 1.345 ;
        RECT 2.06 0.48 2.18 0.54 ;
        RECT 2.435 0.815 2.495 1.345 ;
        RECT 2.47 0.48 2.59 0.555 ;
        RECT 2.845 0.815 2.905 1.345 ;
        RECT 2.91 0.435 2.97 0.555 ;
        RECT 3.06 0.495 3.14 0.875 ;
        RECT 2.025 0.815 3.315 0.875 ;
        RECT 3.255 0.815 3.315 1.345 ;
        RECT 2.135 0.495 3.335 0.555 ;
        RECT 3.29 0.48 3.41 0.54 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.27 0.865 0.33 1.23 ;
        RECT 1.635 0.775 1.695 1.23 ;
        RECT 0.27 1.17 1.695 1.23 ;
        RECT 1.635 0.775 1.74 0.895 ;
        RECT 1.635 0.815 1.765 0.895 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 1.07 ;
        RECT 0.46 0.92 0.58 1.07 ;
        RECT 1.475 0.9 1.535 1.07 ;
        RECT 0.46 1.01 1.535 1.07 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.625 1.365 0.705 ;
        RECT 1.305 0.625 1.365 0.91 ;
        RECT 0.68 0.85 1.365 0.91 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 0.625 0.965 0.75 ;
        RECT 0.68 0.67 1.135 0.75 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.6 0.06 ;
    END
  END VSS
END OR4X8

MACRO DFFSHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX1 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.06 0.6 0.3 0.66 ;
        RECT 0.24 0.54 0.3 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.465 0.805 4.715 0.885 ;
        RECT 4.635 0.805 4.715 1.085 ;
        RECT 4.635 1.005 4.765 1.085 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.225 0.795 4.365 1.085 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.36 1.32 0.97 ;
        RECT 0.965 0.91 1.32 0.97 ;
        RECT 1.26 0.6 1.34 0.73 ;
        RECT 1.26 0.36 2.62 0.42 ;
        RECT 2.56 0.36 2.62 0.74 ;
        RECT 2.56 0.68 2.84 0.74 ;
        RECT 2.78 0.68 2.84 0.8 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END DFFSHQX1

MACRO SDFFSHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX1 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.57 0.56 1.02 ;
        RECT 0.48 0.57 0.6 0.65 ;
        RECT 0.48 0.79 0.74 0.87 ;
        RECT 0.66 0.79 0.74 0.92 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.25 0.635 6.16 0.715 ;
        RECT 6.06 0.6 6.14 0.73 ;
        RECT 6.06 0.61 6.16 0.73 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.535 0.815 5.905 0.935 ;
        RECT 5.825 0.815 5.905 1.025 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.56 0.625 4.83 0.775 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.385 0.875 4.66 1.01 ;
        RECT 4.385 0.875 4.83 0.955 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.98 1.14 1.11 ;
        RECT 1.08 0.875 1.14 1.295 ;
        RECT 1.08 1.235 1.565 1.295 ;
        RECT 1.505 1.22 2.05 1.28 ;
        RECT 1.99 1.12 2.05 1.28 ;
        RECT 2.385 0.915 2.445 1.18 ;
        RECT 1.99 1.12 2.445 1.18 ;
        RECT 2.385 0.915 2.505 0.975 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END SDFFSHQX1

MACRO SDFFSHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX4 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.025 0.655 6.94 0.715 ;
        RECT 6.86 0.6 6.94 0.73 ;
        RECT 6.86 0.645 6.98 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.315 0.815 6.395 0.95 ;
        RECT 6.315 0.815 6.76 0.895 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.235 0.625 5.545 0.705 ;
        RECT 5.465 0.625 5.545 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.015 0.605 5.135 0.685 ;
        RECT 5.035 0.605 5.135 0.895 ;
        RECT 5.035 0.815 5.305 0.895 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.48 0.835 1.54 1.305 ;
        RECT 1.46 1.17 1.54 1.3 ;
        RECT 1.48 0.835 1.67 0.895 ;
        RECT 1.48 1.245 2 1.305 ;
        RECT 1.94 1.205 3.065 1.265 ;
        RECT 3.005 1 3.065 1.265 ;
        RECT 3.005 1 3.125 1.06 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.54 0.495 1.355 ;
        RECT 0.435 0.6 0.54 0.73 ;
        RECT 0.435 0.645 0.86 0.705 ;
        RECT 0.8 0.6 0.86 0.97 ;
        RECT 0.845 0.54 0.905 0.66 ;
        RECT 0.845 0.91 0.905 1.355 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.2 0.06 ;
    END
  END VSS
END SDFFSHQX4

MACRO TLATNTSCAX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX2 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.41 3.34 1.29 ;
        RECT 3.26 0.41 3.36 0.53 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.74 0.95 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.45 0.54 0.95 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.10 0.51 0.2 0.95 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END TLATNTSCAX2

MACRO XNOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.5 0.32 1.465 ;
        RECT 0.26 0.98 0.335 1.465 ;
        RECT 0.26 0.98 0.34 1.135 ;
        RECT 0.245 0.5 0.365 0.56 ;
        RECT 0.26 1.075 0.7 1.135 ;
        RECT 0.64 0.39 0.7 0.61 ;
        RECT 0.26 0.55 0.7 0.61 ;
        RECT 0.64 1.075 0.7 1.405 ;
        RECT 0.685 0.33 0.745 0.45 ;
        RECT 0.685 1.345 0.745 1.465 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.425 0.65 1.485 0.825 ;
        RECT 1.805 0.645 1.865 0.825 ;
        RECT 1.715 0.765 1.835 0.91 ;
        RECT 1.425 0.765 1.865 0.825 ;
        RECT 1.835 0.625 2.08 0.705 ;
        RECT 2.02 0.625 2.08 0.745 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.96 0.71 1.165 1.085 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END XNOR2X4

MACRO DFFSX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX2 0 0 ;
  SIZE 6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.57 5.34 1.29 ;
        RECT 5.23 0.57 5.35 0.65 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.62 0.55 4.74 0.63 ;
        RECT 4.66 0.55 4.74 1.29 ;
    END
  END Q
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 0.75 3.54 1.25 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6 0.06 ;
    END
  END VSS
END DFFSX2

MACRO DFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.6 3.74 0.73 ;
        RECT 3.66 0.645 3.9 0.705 ;
        RECT 3.84 0.53 3.9 1.29 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.53 3.34 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.53 2.94 1.03 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 0.935 0.365 1.275 ;
        RECT 0.235 1.195 0.365 1.275 ;
        RECT 0.37 0.895 0.45 1.015 ;
        RECT 0.285 0.935 0.45 1.015 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END DFFX2

MACRO SEDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFX2 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.1 0.4 6.18 1.11 ;
        RECT 6.06 0.98 6.18 1.11 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.28 0.54 0.34 1.29 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.675 0.585 6.735 1.085 ;
        RECT 6.675 0.585 6.795 0.65 ;
        RECT 6.675 0.585 7.485 0.645 ;
        RECT 7.425 0.625 7.565 0.705 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.895 0.745 7.165 0.895 ;
        RECT 6.895 0.745 7.325 0.825 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.635 0.61 5.765 0.98 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.235 0.815 4.365 0.895 ;
        RECT 4.285 0.815 4.365 1.265 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.755 3.94 0.92 ;
        RECT 3.86 0.84 4.135 0.92 ;
        RECT 4.055 0.84 4.135 1.06 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.8 0.06 ;
    END
  END VSS
END SEDFFX2

MACRO ADDFHXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHXL 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.085 0.51 4.145 1.405 ;
        RECT 4.085 0.6 4.34 0.73 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.6 0.14 0.98 ;
        RECT 0.08 0.92 0.405 0.98 ;
        RECT 0.345 0.465 0.405 0.66 ;
        RECT 0.06 0.6 0.405 0.66 ;
        RECT 0.345 0.92 0.405 1.21 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.625 1.025 2.74 1.045 ;
        RECT 1.07 0.965 1.765 1.025 ;
        RECT 1.705 1.025 2.74 1.085 ;
        RECT 2.68 0.965 3.535 1.025 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.905 0.805 0.965 0.925 ;
        RECT 0.905 0.805 1.915 0.865 ;
        RECT 0.905 0.825 1.985 0.865 ;
        RECT 1.865 0.865 2.58 0.925 ;
        RECT 2.52 0.805 3.765 0.865 ;
        RECT 3.635 0.805 3.765 0.895 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.53 0.625 1.765 0.705 ;
        RECT 2.11 0.645 2.17 0.765 ;
        RECT 1.53 0.645 3.235 0.705 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END ADDFHXL

MACRO OAI221X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X2 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 1.155 0.72 1.275 ;
        RECT 1.68 1.155 1.74 1.275 ;
        RECT 2.34 1.155 2.4 1.405 ;
        RECT 2.44 0.475 2.5 1.215 ;
        RECT 0.66 1.155 2.5 1.215 ;
        RECT 2.44 0.79 2.54 0.92 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.22 0.86 0.34 0.92 ;
        RECT 0.28 0.79 0.34 1.055 ;
        RECT 0.94 0.845 1 1.055 ;
        RECT 0.28 0.995 1 1.055 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.4 0.845 1.46 1.055 ;
        RECT 2.06 0.79 2.14 1.055 ;
        RECT 1.4 0.995 2.14 1.055 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.715 0.715 0.795 ;
        RECT 0.635 0.715 0.715 0.895 ;
        RECT 0.635 0.815 0.84 0.895 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.685 0.715 1.765 0.895 ;
        RECT 1.56 0.815 1.765 0.895 ;
        RECT 1.685 0.715 1.96 0.795 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.555 2.34 1.055 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END OAI221X2

MACRO SEDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX2 0 0 ;
  SIZE 7.0 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.495 3.14 1.025 ;
        RECT 3.06 0.495 3.185 0.575 ;
        RECT 3.06 0.945 3.265 1.025 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.48 0.67 6.56 0.96 ;
        RECT 6.48 0.79 6.77 0.96 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.705 2.96 0.92 ;
        RECT 2.88 0.705 2.96 1.185 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.625 0.625 1.775 0.895 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.585 0.74 1.085 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.365 0.705 ;
        RECT 0.5 0.425 0.56 0.685 ;
        RECT 0.235 0.625 0.56 0.685 ;
        RECT 0.5 0.425 0.96 0.485 ;
        RECT 0.9 0.425 0.96 0.655 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.8 0.06 ;
    END
  END VSS
END SEDFFHQX2

MACRO SDFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRX1 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.41 1 0.54 ;
        RECT 0.94 0.41 1 1.33 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.29 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.06 0.43 6.14 0.735 ;
        RECT 5.865 0.6 6.14 0.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.62 0.46 5.7 0.895 ;
        RECT 5.62 0.815 5.765 0.895 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.19 0.625 5.365 0.875 ;
        RECT 5.19 0.625 5.52 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.86 0.625 3.94 0.92 ;
        RECT 3.86 0.785 4.145 0.92 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.285 0.77 1.365 1.085 ;
        RECT 1.1 1.005 1.365 1.085 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END SDFFTRX1

MACRO AND4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.305 0.295 1.365 0.415 ;
        RECT 1.305 0.815 1.365 1.335 ;
        RECT 1.305 0.355 1.46 0.415 ;
        RECT 1.4 0.355 1.46 0.875 ;
        RECT 1.305 0.815 1.46 0.875 ;
        RECT 1.4 0.6 1.54 0.73 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.675 1.08 0.92 ;
        RECT 1.06 0.775 1.14 1.115 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 1.1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.035 0.625 0.36 0.995 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END AND4X2

MACRO OAI22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.98 0.54 1.11 ;
        RECT 0.48 0.64 0.54 1.235 ;
        RECT 0.635 0.45 0.695 0.7 ;
        RECT 0.48 0.64 0.695 0.7 ;
        RECT 0.735 0.39 0.795 0.51 ;
        RECT 0.635 0.45 0.795 0.51 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 1.05 ;
        RECT 0.29 0.58 0.37 0.92 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 1.1 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.61 0.94 1.11 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.8 0.74 1.3 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OAI22XL

MACRO DFFSHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.285 0.445 5.365 0.895 ;
        RECT 5.235 0.815 5.365 0.895 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.385 0.715 4.465 0.895 ;
        RECT 4.385 0.815 4.785 0.895 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.355 1.92 0.925 ;
        RECT 1.445 0.865 1.92 0.925 ;
        RECT 1.86 0.6 1.94 0.73 ;
        RECT 1.86 0.355 2.81 0.415 ;
        RECT 2.75 0.355 2.81 0.575 ;
        RECT 2.75 0.515 3.075 0.575 ;
        RECT 3.015 0.515 3.075 0.7 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.365 0.73 ;
        RECT 0.305 0.54 0.365 1.465 ;
        RECT 0.26 0.67 0.775 0.73 ;
        RECT 0.715 0.54 0.775 1.465 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.6 0.06 ;
    END
  END VSS
END DFFSHQX4

MACRO NOR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2XL 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.37 0.32 0.49 ;
        RECT 0.26 0.43 0.57 0.49 ;
        RECT 0.51 0.43 0.57 1.145 ;
        RECT 0.46 0.98 0.57 1.145 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.16 0.54 ;
        RECT 0.08 0.41 0.16 0.89 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 1.02 ;
        RECT 0.33 0.59 0.41 0.87 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.6 0.06 ;
    END
  END VSS
END NOR2XL

MACRO XNOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X2 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.54 0.54 1.12 ;
        RECT 0.42 1.04 0.54 1.12 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.59 0.815 2.09 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.685 0.905 0.895 ;
        RECT 0.64 0.815 1.01 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END XNOR2X2

MACRO INVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1 0 0 ;
  SIZE 0.40 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 0.72 0.335 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.72 0.155 0.8 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.40 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.40 0.06 ;
    END
  END VSS
END INVX1

MACRO NAND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X8 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 0.995 0.355 1.44 ;
        RECT 0.705 1.05 0.765 1.44 ;
        RECT 1.115 1.05 1.175 1.44 ;
        RECT 1.525 1.05 1.585 1.44 ;
        RECT 1.935 1.05 1.995 1.44 ;
        RECT 2.345 1.05 2.405 1.44 ;
        RECT 2.755 1.05 2.815 1.44 ;
        RECT 0.47 0.545 3.14 0.605 ;
        RECT 3.06 0.98 3.14 1.11 ;
        RECT 3.08 0.545 3.14 1.11 ;
        RECT 0.295 1.05 3.14 1.11 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.535 0.865 0.81 0.925 ;
        RECT 1.43 0.865 1.55 0.95 ;
        RECT 2.045 0.865 2.165 0.95 ;
        RECT 2.635 0.815 2.765 0.95 ;
        RECT 0.75 0.89 2.765 0.95 ;
        RECT 2.635 0.815 2.875 0.875 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.365 0.79 ;
        RECT 0.91 0.705 1.03 0.79 ;
        RECT 1.775 0.705 1.895 0.79 ;
        RECT 0.235 0.705 2.325 0.765 ;
        RECT 2.265 0.73 2.51 0.79 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END NAND2X8

MACRO SDFFQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.515 0.645 4.575 0.985 ;
        RECT 4.455 0.925 4.575 0.985 ;
        RECT 5.035 0.625 5.165 0.705 ;
        RECT 4.515 0.645 5.165 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.835 0.805 4.94 1.015 ;
        RECT 4.835 0.805 5.205 0.895 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.005 0.755 4.165 0.895 ;
        RECT 4.085 0.755 4.165 0.985 ;
        RECT 4.005 0.755 4.355 0.875 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.65 0.31 0.97 ;
        RECT 0.26 0.5 0.34 0.73 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.57 0.73 ;
        RECT 0.51 0.57 0.57 1.29 ;
        RECT 0.48 0.57 0.6 0.66 ;
        RECT 0.46 0.6 0.935 0.66 ;
        RECT 0.875 0.57 0.935 0.945 ;
        RECT 0.92 0.885 0.98 1.29 ;
        RECT 0.875 0.57 1.07 0.63 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END SDFFQX4

MACRO SDFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFXL 0 0 ;
  SIZE 5.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.54 0.94 1.21 ;
        RECT 1.035 0.5 1.115 0.62 ;
        RECT 0.86 0.54 1.115 0.62 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.305 0.635 ;
        RECT 0.225 0.41 0.305 1.02 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.78 0.835 4.84 1.01 ;
        RECT 4.8 0.585 4.86 0.895 ;
        RECT 4.8 0.585 5.105 0.705 ;
        RECT 5.325 0.585 5.385 0.705 ;
        RECT 4.8 0.625 5.385 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.96 0.805 5.385 0.895 ;
        RECT 5.235 0.805 5.385 0.96 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.68 4.34 0.96 ;
        RECT 4.26 0.785 4.52 0.92 ;
        RECT 4.44 0.785 4.52 0.96 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.285 0.88 1.365 1.085 ;
        RECT 1.04 1.005 1.365 1.085 ;
        RECT 1.285 0.88 1.415 0.96 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.8 0.06 ;
    END
  END VSS
END SDFFXL

MACRO CLKBUFX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX20 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.355 0.13 1.36 ;
        RECT 0.06 0.595 0.14 0.975 ;
        RECT 0.48 0.355 0.54 0.655 ;
        RECT 0.48 0.915 0.54 1.36 ;
        RECT 0.89 0.355 0.95 0.655 ;
        RECT 0.89 0.915 0.95 1.36 ;
        RECT 1.3 0.355 1.36 0.655 ;
        RECT 1.3 0.915 1.36 1.36 ;
        RECT 1.71 0.355 1.77 0.655 ;
        RECT 1.71 0.915 1.77 1.36 ;
        RECT 2.12 0.355 2.18 0.655 ;
        RECT 2.12 0.915 2.18 1.36 ;
        RECT 2.53 0.355 2.59 0.655 ;
        RECT 2.53 0.915 2.59 1.36 ;
        RECT 2.94 0.355 3 0.655 ;
        RECT 2.94 0.915 3 1.36 ;
        RECT 0.06 0.915 3.41 0.975 ;
        RECT 3.35 0.355 3.41 0.655 ;
        RECT 0.06 0.595 3.41 0.655 ;
        RECT 3.35 0.915 3.41 1.36 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.875 0.815 4.375 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END CLKBUFX20

MACRO OAI2BB2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 1.005 1.565 1.085 ;
        RECT 1.64 1.025 1.7 1.455 ;
        RECT 1.435 1.025 2.135 1.085 ;
        RECT 2.075 0.58 2.135 1.265 ;
        RECT 2.28 0.4 2.34 0.64 ;
        RECT 2.28 0.4 2.4 0.46 ;
        RECT 2.075 1.205 2.53 1.265 ;
        RECT 2.47 1.205 2.53 1.325 ;
        RECT 2.675 0.4 2.735 0.64 ;
        RECT 2.075 0.58 2.735 0.64 ;
        RECT 2.675 0.4 2.81 0.46 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.465 0.815 2.84 0.895 ;
        RECT 2.635 0.74 2.84 0.945 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.775 2.295 1.105 ;
        RECT 2.235 0.815 2.365 0.895 ;
        RECT 2.94 0.87 3 1.105 ;
        RECT 2.235 1.045 3 1.105 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 0.625 0.725 0.895 ;
        RECT 0.415 0.815 0.725 0.895 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.315 0.895 ;
        RECT 0.235 0.625 0.545 0.705 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END OAI2BB2X2

MACRO FILL32
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL32 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END FILL32

MACRO OAI33X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.785 1.21 0.845 1.46 ;
        RECT 0.99 0.37 1.05 0.51 ;
        RECT 1.4 0.37 1.5 0.51 ;
        RECT 0.99 0.45 1.5 0.51 ;
        RECT 1.44 0.37 1.5 1.27 ;
        RECT 1.44 0.98 1.54 1.27 ;
        RECT 0.785 1.21 1.54 1.27 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.61 0.94 1.11 ;
    END
  END B2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END A0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.61 0.74 1.11 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.61 1.14 1.11 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.61 1.34 1.11 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END OAI33X1

MACRO SDFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRX4 0 0 ;
  SIZE 7.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.27 0.485 6.34 1.29 ;
        RECT 6.26 0.79 6.34 1.29 ;
        RECT 6.26 0.9 6.75 0.96 ;
        RECT 6.69 0.9 6.75 1.29 ;
        RECT 6.27 0.485 6.86 0.545 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.46 0.79 5.52 1.29 ;
        RECT 5.48 0.485 5.54 0.96 ;
        RECT 5.46 0.9 5.93 0.96 ;
        RECT 5.33 0.485 5.92 0.545 ;
        RECT 5.87 0.9 5.93 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.24 0.525 2.32 0.87 ;
        RECT 2.26 0.79 2.34 1.005 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.995 0.525 2.075 0.87 ;
        RECT 2.06 0.79 2.14 0.96 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.945 0.625 1.165 0.91 ;
        RECT 0.87 0.815 1.165 0.91 ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.625 0.77 0.745 ;
        RECT 0.69 0.625 0.77 1.07 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 0.92 ;
        RECT 0.295 0.655 0.375 0.87 ;
        RECT 0.06 0.79 0.375 0.87 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.6 0.06 ;
    END
  END VSS
END SDFFTRX4

MACRO NOR2BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BXL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.48 0.14 1.3 ;
        RECT 0.06 1.17 0.14 1.3 ;
        RECT 0.06 1.24 0.29 1.3 ;
        RECT 0.23 1.24 0.29 1.36 ;
        RECT 0.335 0.285 0.395 0.54 ;
        RECT 0.08 0.48 0.395 0.54 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.98 0.54 1.11 ;
        RECT 0.565 0.715 0.645 1.06 ;
        RECT 0.46 0.98 0.645 1.06 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.64 0.34 1.14 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END NOR2BXL

MACRO MXI2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.485 0.72 1.365 ;
        RECT 0.66 0.79 0.74 0.92 ;
        RECT 0.66 0.485 0.855 0.545 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.5 0.325 0.56 0.935 ;
        RECT 0.5 0.325 1.015 0.385 ;
        RECT 0.955 0.325 1.015 0.705 ;
        RECT 0.83 0.645 1.365 0.705 ;
        RECT 1.16 0.625 1.365 0.715 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.815 1.14 0.985 ;
        RECT 1 0.815 1.41 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.535 0.34 1.035 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END MXI2X1

MACRO NOR4BBX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.465 1.345 0.525 1.465 ;
        RECT 0.595 0.465 0.715 0.525 ;
        RECT 0.665 0.485 1.12 0.545 ;
        RECT 1.06 0.425 1.12 1.405 ;
        RECT 0.465 1.345 1.12 1.405 ;
        RECT 1.06 0.98 1.14 1.11 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.845 0.54 1.245 ;
        RECT 0.495 0.805 0.6 0.925 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.805 0.78 1.06 ;
        RECT 0.7 0.98 0.94 1.06 ;
        RECT 0.86 0.98 0.94 1.145 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.815 1.565 1.07 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.08 0.46 0.16 0.89 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END NOR4BBX1

MACRO CLKINVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX2 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.52 0.54 1.29 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.76 ;
        RECT 0.06 0.68 0.36 0.76 ;
        RECT 0.28 0.6 0.36 0.8 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.8 0.06 ;
    END
  END VSS
END CLKINVX2

MACRO SDFFQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.365 0.73 ;
        RECT 0.305 0.37 0.365 1.29 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.75 0.785 3.81 0.96 ;
        RECT 3.775 0.645 3.835 0.845 ;
        RECT 4.035 0.625 4.165 0.705 ;
        RECT 3.775 0.645 4.48 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.2 0.805 4.61 0.895 ;
        RECT 4.435 0.805 4.61 0.975 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.625 3.34 0.975 ;
        RECT 3.26 0.79 3.49 0.92 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.61 0.74 1.11 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END SDFFQX2

MACRO AOI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 0.37 0.74 1.11 ;
        RECT 0.66 0.98 0.74 1.11 ;
        RECT 0.66 1.05 0.995 1.11 ;
        RECT 0.935 1.05 0.995 1.19 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.45 1.14 0.95 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.41 0.94 0.91 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.54 0.35 ;
        RECT 0.48 0.27 0.56 0.7 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END AOI22X1

MACRO TLATNTSCAX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX20 0 0 ;
  SIZE 8.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.355 5.32 1.36 ;
        RECT 5.26 0.76 5.34 1.36 ;
        RECT 5.67 0.355 5.73 1.36 ;
        RECT 6.035 0.6 6.095 0.82 ;
        RECT 6.08 0.355 6.14 0.66 ;
        RECT 6.08 0.76 6.14 1.36 ;
        RECT 6.49 0.355 6.55 1.36 ;
        RECT 6.9 0.355 6.96 1.36 ;
        RECT 7.31 0.355 7.37 1.36 ;
        RECT 7.72 0.355 7.78 1.36 ;
        RECT 8.13 0.355 8.19 1.36 ;
        RECT 5.26 0.76 8.6 0.82 ;
        RECT 8.495 0.6 8.555 0.82 ;
        RECT 8.54 0.355 8.6 0.66 ;
        RECT 8.54 0.76 8.6 1.355 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.74 0.67 0.965 0.895 ;
        RECT 0.695 0.815 1.05 0.895 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 0.955 ;
        RECT 0.515 0.51 0.595 0.87 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.98 0.14 1.14 ;
        RECT 0.12 0.7 0.2 1.06 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 8.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 8.8 0.06 ;
    END
  END VSS
END TLATNTSCAX20

MACRO AO21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.405 1.14 0.99 ;
        RECT 1.06 0.91 1.295 0.99 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.6 0.16 1.08 ;
        RECT 0.06 0.79 0.16 1.08 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.34 0.92 ;
        RECT 0.44 0.6 0.52 0.87 ;
        RECT 0.26 0.79 0.52 0.87 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.62 0.73 0.74 0.81 ;
        RECT 0.66 0.73 0.74 1.19 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END AO21XL

MACRO OAI32XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 1.005 1.165 1.085 ;
        RECT 1.105 0.74 1.165 1.235 ;
        RECT 1.24 0.415 1.3 0.8 ;
        RECT 1.105 0.74 1.3 0.8 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.56 0.92 ;
        RECT 0.48 0.79 0.56 1.27 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 0.9 1.345 1.11 ;
        RECT 1.46 0.935 1.54 1.11 ;
        RECT 1.265 1.03 1.54 1.11 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.74 0.74 0.975 ;
        RECT 0.66 0.74 1.005 0.82 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.425 0.655 1.505 0.8 ;
        RECT 1.425 0.72 1.74 0.8 ;
        RECT 1.66 0.72 1.74 0.92 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OAI32XL

MACRO NOR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.505 0.465 0.76 ;
        RECT 0.405 0.7 0.92 0.76 ;
        RECT 0.84 1.115 0.9 1.235 ;
        RECT 0.86 0.505 0.92 1.175 ;
        RECT 0.86 0.505 0.94 0.73 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.935 0.74 1.355 ;
        RECT 0.665 0.86 0.745 1.015 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.03 0.86 0.11 1.11 ;
        RECT 0.03 0.955 0.36 1.11 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.945 0.54 1.445 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END NOR3XL

MACRO EDFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRXL 0 0 ;
  SIZE 6.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.52 0.94 1.02 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.285 0.73 ;
        RECT 0.205 0.54 0.285 1.02 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.23 0.735 6.435 0.855 ;
        RECT 6.26 0.735 6.435 1.11 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.405 0.765 5.965 0.845 ;
        RECT 5.835 0.765 5.965 0.895 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.29 0.85 4.54 0.93 ;
        RECT 4.46 0.85 4.54 1.18 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.545 1.14 0.77 ;
        RECT 1.085 0.69 1.165 1.02 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.8 0.06 ;
    END
  END VSS
END EDFFTRXL

MACRO MX4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X2 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.6 1.74 1.04 ;
        RECT 1.6 0.96 1.74 1.04 ;
        RECT 1.67 0.425 1.75 0.68 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.04 0.59 4.1 0.71 ;
        RECT 4.04 0.59 4.72 0.65 ;
        RECT 4.66 0.59 4.72 0.92 ;
        RECT 4.66 0.79 4.74 0.92 ;
    END
  END S0
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.2 0.75 4.28 0.97 ;
        RECT 4.2 0.75 4.56 0.895 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.98 3.34 1.28 ;
        RECT 3.32 0.84 3.4 1.06 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.92 0.84 3 1.28 ;
        RECT 2.86 0.965 3 1.28 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.79 1.94 0.92 ;
        RECT 2.095 0.655 2.175 0.87 ;
        RECT 1.86 0.79 2.175 0.87 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.17 0.62 1.27 0.87 ;
        RECT 1.26 0.46 1.34 0.73 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END MX4X2

MACRO NAND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X6 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 1.015 0.465 1.345 ;
        RECT 0.64 0.435 0.7 0.555 ;
        RECT 0.815 1.015 0.875 1.345 ;
        RECT 1.235 1.015 1.295 1.345 ;
        RECT 1.54 0.435 1.6 0.555 ;
        RECT 1.645 1.015 1.705 1.345 ;
        RECT 2.055 1.015 2.115 1.345 ;
        RECT 2.16 0.435 2.22 0.555 ;
        RECT 0.405 1.015 2.76 1.075 ;
        RECT 2.465 1.015 2.525 1.345 ;
        RECT 0.64 0.495 2.76 0.555 ;
        RECT 2.66 0.98 2.74 1.11 ;
        RECT 2.7 0.495 2.76 1.085 ;
        RECT 2.465 1.015 2.76 1.085 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.71 0.815 0.975 0.875 ;
        RECT 1.445 0.815 1.565 0.915 ;
        RECT 0.915 0.855 2.085 0.915 ;
        RECT 2.035 0.815 2.185 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.54 0.755 ;
        RECT 0.345 0.695 0.54 0.755 ;
        RECT 1.075 0.655 1.195 0.755 ;
        RECT 1.755 0.655 1.875 0.745 ;
        RECT 0.46 0.655 2.6 0.715 ;
        RECT 2.54 0.655 2.6 0.88 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END NAND2X6

MACRO AOI21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.405 0.7 0.63 ;
        RECT 0.64 0.57 0.92 0.63 ;
        RECT 0.84 1.235 0.9 1.355 ;
        RECT 0.86 0.57 0.92 1.295 ;
        RECT 0.86 0.6 0.94 0.73 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.88 ;
        RECT 0.06 0.61 0.36 0.69 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.54 0.72 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.73 0.74 1.23 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1 0.06 ;
    END
  END VSS
END AOI21XL

MACRO NAND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X4 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 0.995 0.4 1.345 ;
        RECT 0.63 0.475 0.75 0.535 ;
        RECT 0.75 0.995 0.81 1.345 ;
        RECT 1.16 0.995 1.22 1.345 ;
        RECT 1.25 0.475 1.37 0.555 ;
        RECT 1.57 0.995 1.63 1.345 ;
        RECT 0.7 0.495 1.765 0.555 ;
        RECT 1.635 0.815 1.765 0.895 ;
        RECT 1.705 0.495 1.765 1.055 ;
        RECT 0.34 0.995 1.765 1.055 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 0.815 1.295 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.365 0.715 ;
        RECT 0.235 0.655 1.605 0.715 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END NAND2X4

MACRO NOR4BBX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 0.36 1.315 0.48 ;
        RECT 1.665 0.36 1.725 0.48 ;
        RECT 2.075 0.36 2.135 0.48 ;
        RECT 2.485 0.36 2.545 0.48 ;
        RECT 2.925 0.36 2.985 0.48 ;
        RECT 3.335 0.36 3.395 0.48 ;
        RECT 3.775 0.36 3.835 0.48 ;
        RECT 1.255 0.42 3.9 0.48 ;
        RECT 3.84 0.42 3.9 1.3 ;
        RECT 3.84 0.98 3.94 1.11 ;
        RECT 4.185 0.37 4.245 0.51 ;
        RECT 3.84 0.45 4.245 0.51 ;
        RECT 3.84 0.98 4.31 1.04 ;
        RECT 4.25 0.98 4.31 1.3 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.61 3.74 1.11 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.58 2.94 1.08 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.76 0.54 1.26 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.76 0.34 1.26 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END NOR4BBX4

MACRO SDFFSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRXL 0 0 ;
  SIZE 7.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 0.73 ;
        RECT 0.88 0.55 0.94 1.255 ;
        RECT 0.935 0.515 0.995 0.635 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 0.53 0.26 0.73 ;
        RECT 0.06 0.6 0.26 0.73 ;
        RECT 0.18 0.53 0.26 0.99 ;
        RECT 0.23 0.405 0.31 0.62 ;
        RECT 0.23 0.9 0.31 1.02 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.715 0.655 6.775 1 ;
        RECT 6.895 0.595 6.955 0.715 ;
        RECT 7.275 0.595 7.335 0.715 ;
        RECT 7.235 0.625 7.365 0.715 ;
        RECT 6.715 0.655 7.365 0.715 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.035 0.815 7.275 0.985 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.235 0.815 6.455 0.895 ;
        RECT 6.375 0.815 6.455 1.175 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.775 1.005 6.275 1.085 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.815 2.365 0.895 ;
        RECT 2.1 0.835 2.365 0.895 ;
        RECT 2.305 0.815 2.365 1.01 ;
        RECT 2.305 0.95 3.15 1.01 ;
        RECT 3.09 0.95 3.15 1.24 ;
        RECT 3.09 1.18 4.06 1.24 ;
        RECT 4 1.18 4.06 1.4 ;
        RECT 4 1.34 4.485 1.4 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.04 0.9 1.365 1.085 ;
        RECT 1.245 0.995 1.39 1.13 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.6 0.06 ;
    END
  END VSS
END SDFFSRXL

MACRO OR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.37 1.14 1.3 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.625 0.8 1.04 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.645 0.375 0.92 ;
        RECT 0.295 0.645 0.375 1.11 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.61 0.14 1.11 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OR3X1

MACRO AOI211X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 0.445 0.67 0.505 ;
        RECT 1.06 0.465 1.14 0.73 ;
        RECT 1.08 0.465 1.14 1.005 ;
        RECT 1.195 0.445 1.315 0.525 ;
        RECT 1.08 0.945 1.725 1.005 ;
        RECT 0.62 0.465 1.685 0.525 ;
        RECT 1.665 0.945 1.725 1.225 ;
        RECT 1.635 0.445 1.755 0.505 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.525 0.805 0.895 0.915 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.905 0.705 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.625 1.6 0.705 ;
        RECT 1.435 0.625 1.6 0.845 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.7 0.625 1.965 0.795 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END AOI211X2

MACRO BUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX6 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.57 1.54 1.07 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.35 0.13 1.37 ;
        RECT 0.06 0.79 0.14 0.975 ;
        RECT 0.48 0.35 0.54 0.655 ;
        RECT 0.48 0.915 0.54 1.37 ;
        RECT 0.06 0.915 0.95 0.975 ;
        RECT 0.89 0.35 0.95 0.655 ;
        RECT 0.06 0.595 0.95 0.655 ;
        RECT 0.89 0.915 0.95 1.37 ;
    END
  END Y
END BUFX6

MACRO NOR3BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BXL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.47 0.14 1.29 ;
        RECT 0.14 0.275 0.2 0.53 ;
        RECT 0.08 1.23 0.275 1.29 ;
        RECT 0.215 1.23 0.275 1.35 ;
        RECT 0.505 0.305 0.565 0.53 ;
        RECT 0.08 0.47 0.565 0.53 ;
        RECT 0.505 0.305 0.64 0.365 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.765 0.775 0.845 1.13 ;
        RECT 0.825 0.75 0.905 0.895 ;
        RECT 0.765 0.775 0.965 0.895 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.63 0.54 1.13 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.63 0.34 1.13 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END NOR3BXL

MACRO MXI3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3X1 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.54 3.74 1.29 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.235 0.62 3.315 0.86 ;
        RECT 3.06 0.62 3.4 0.74 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.8 2.355 0.99 ;
        RECT 2.235 0.815 2.365 0.99 ;
        RECT 2.235 0.91 2.765 0.99 ;
    END
  END S1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.42 0.84 1.5 1.085 ;
        RECT 1.42 1.005 1.755 1.085 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.37 0.775 0.565 0.905 ;
        RECT 0.37 0.775 0.82 0.855 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.19 0.895 0.27 1.085 ;
        RECT 0.92 0.93 1 1.085 ;
        RECT 0.19 1.005 1 1.085 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.8 0.06 ;
    END
  END VSS
END MXI3X1

MACRO NAND2BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX2 0 0 ;
  SIZE 1.20 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.075 0.55 0.155 0.635 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.775 1.115 0.935 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.075 0.955 0.155 1.035 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.20 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.20 0.06 ;
    END
  END VSS
END NAND2BX2

MACRO AOI32X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.85 0.505 0.91 1.085 ;
        RECT 0.85 1.005 1.165 1.085 ;
        RECT 1.105 1.005 1.165 1.305 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.48 0.48 0.56 0.89 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.625 1.315 0.85 ;
        RECT 1.01 0.77 1.315 0.85 ;
        RECT 1.235 0.625 1.365 0.705 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.41 0.74 0.54 ;
        RECT 0.67 0.46 0.75 0.9 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 0.65 1.545 0.905 ;
        RECT 1.66 0.6 1.74 0.73 ;
        RECT 1.465 0.65 1.74 0.73 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.585 0.34 1.085 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END AOI32X1

MACRO OAI2BB1XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 0.54 ;
        RECT 0.08 0.3 0.14 0.68 ;
        RECT 0.08 0.62 0.36 0.68 ;
        RECT 0.28 0.24 0.34 0.36 ;
        RECT 0.08 0.3 0.34 0.36 ;
        RECT 0.3 0.62 0.36 1.28 ;
        RECT 0.3 1.22 0.47 1.28 ;
        RECT 0.41 1.22 0.47 1.34 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.62 0.54 1.12 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.62 0.74 1.12 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.61 1.14 1.11 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END OAI2BB1XL

MACRO AO22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.25 0.405 1.33 0.68 ;
        RECT 1.26 0.6 1.34 0.99 ;
        RECT 1.26 0.91 1.51 0.99 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.79 1.14 0.87 ;
        RECT 1.06 0.79 1.14 1.23 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.595 0.74 1.095 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.23 0.54 0.73 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END AO22XL

MACRO NAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X2 0 0 ;
  SIZE 1.00 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.87 0.76 0.95 0.84 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.62 0.57 0.72 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.065 0.8 0.15 0.98 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.00 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.00 0.06 ;
    END
  END VSS
END NAND2X2

MACRO NOR4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.35 0.29 0.41 0.545 ;
        RECT 0.79 0.29 0.85 0.545 ;
        RECT 0.35 0.485 1.14 0.545 ;
        RECT 1.08 0.485 1.14 1.11 ;
        RECT 1.04 0.98 1.14 1.11 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.645 0.36 0.895 ;
        RECT 0.03 0.815 0.36 0.895 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.73 0.54 1.23 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.645 0.74 1.145 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.65 0.94 1.11 ;
        RECT 0.86 0.65 0.98 0.73 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END NOR4XL

MACRO MX3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3XL 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.16 0.54 ;
        RECT 0.1 0.41 0.16 1.29 ;
        RECT 0.04 1.23 0.16 1.29 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.965 0.79 2.045 0.91 ;
        RECT 2.025 0.83 2.105 1.165 ;
        RECT 2.46 0.98 2.54 1.165 ;
        RECT 2.025 1.085 2.54 1.165 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.74 2.34 0.985 ;
        RECT 2.205 0.74 2.54 0.82 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.575 1.54 0.775 ;
        RECT 1.465 0.6 1.545 1.07 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.575 1.34 1.07 ;
        RECT 1.255 0.95 1.34 1.07 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.765 0.34 1.195 ;
        RECT 0.26 0.765 0.41 0.885 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END MX3XL

MACRO CLKINVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX8 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.995 0.385 1.345 ;
        RECT 0.295 0.57 0.415 0.63 ;
        RECT 0.735 0.995 0.795 1.345 ;
        RECT 0.705 0.57 0.825 0.645 ;
        RECT 0.325 0.995 1.205 1.055 ;
        RECT 1.145 0.525 1.205 0.645 ;
        RECT 1.145 0.96 1.205 1.345 ;
        RECT 1.26 0.585 1.32 1.02 ;
        RECT 1.26 0.585 1.34 0.73 ;
        RECT 1.135 0.96 1.615 1.02 ;
        RECT 0.37 0.585 1.57 0.645 ;
        RECT 1.555 0.96 1.615 1.345 ;
        RECT 1.525 0.57 1.645 0.63 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.77 0.565 0.895 ;
        RECT 0.435 0.77 1.095 0.85 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END CLKINVX8

MACRO NAND4BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.44 0.14 1.26 ;
        RECT 0.06 0.98 0.14 1.26 ;
        RECT 0.205 0.38 0.265 0.5 ;
        RECT 0.08 0.44 0.265 0.5 ;
        RECT 0.36 1.2 0.42 1.48 ;
        RECT 0.06 1.2 0.84 1.26 ;
        RECT 0.78 1.2 0.84 1.48 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.76 1.14 1.26 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.43 0.73 0.92 ;
        RECT 0.65 0.79 0.74 0.92 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 0.92 ;
        RECT 0.47 0.8 0.55 1.1 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END NAND4BX1

MACRO AOI31XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.9 0.54 0.96 0.795 ;
        RECT 0.9 0.735 1.325 0.795 ;
        RECT 1.265 0.735 1.325 1.21 ;
        RECT 1.265 0.79 1.54 0.92 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.79 0.34 0.895 ;
        RECT 0.26 0.79 0.34 1.085 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.93 1.165 1.085 ;
        RECT 1.085 0.93 1.165 1.38 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.645 0.8 0.92 ;
        RECT 0.72 0.645 0.8 1.085 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.79 0.54 0.92 ;
        RECT 0.465 0.425 0.545 0.91 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.6 0.06 ;
    END
  END VSS
END AOI31XL

MACRO DLY1X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY1X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.52 1.74 1.29 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 0.775 0.54 0.895 ;
        RECT 0.46 0.62 0.54 0.94 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END DLY1X1

MACRO OAI21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X4 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.63 1.02 0.69 1.375 ;
        RECT 1.25 1.02 1.31 1.375 ;
        RECT 1.86 1.02 1.92 1.375 ;
        RECT 1.875 0.475 1.935 1.3 ;
        RECT 0.63 1.02 1.935 1.08 ;
        RECT 1.86 1.035 1.94 1.3 ;
        RECT 1.875 0.475 2.05 0.585 ;
        RECT 1.86 1.035 2.33 1.095 ;
        RECT 2.27 1.035 2.33 1.375 ;
        RECT 1.875 0.525 2.385 0.585 ;
        RECT 2.325 0.475 2.46 0.535 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.815 0.68 0.91 ;
        RECT 0.435 0.83 1.265 0.91 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.21 0.66 0.335 0.72 ;
        RECT 0.835 0.655 0.955 0.73 ;
        RECT 0.3 0.655 1.635 0.715 ;
        RECT 1.575 0.655 1.635 0.85 ;
        RECT 1.575 0.79 1.74 0.85 ;
        RECT 1.66 0.79 1.74 0.92 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 0.685 2.115 0.935 ;
        RECT 2.035 0.815 2.365 0.895 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END OAI21X4

MACRO SDFFRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX8 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.78 0.645 6.84 0.915 ;
        RECT 6.78 0.645 7.565 0.705 ;
        RECT 7.345 0.625 7.565 0.715 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.13 0.815 7.365 0.915 ;
        RECT 7.13 0.815 7.61 0.895 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.6 6.34 0.73 ;
        RECT 6.26 0.625 6.52 0.705 ;
        RECT 6.44 0.625 6.52 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.545 0.59 3.655 0.915 ;
        RECT 3.4 0.815 3.655 0.915 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.625 1.965 0.765 ;
        RECT 1.905 0.345 1.965 0.765 ;
        RECT 1.805 0.705 1.965 0.765 ;
        RECT 1.905 0.345 2.45 0.405 ;
        RECT 2.39 0.345 2.45 0.755 ;
        RECT 2.39 0.695 2.545 0.755 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.195 0.67 0.255 1.35 ;
        RECT 0.26 0.54 0.34 0.73 ;
        RECT 0.605 0.67 0.665 1.35 ;
        RECT 0.69 0.54 0.75 0.73 ;
        RECT 1.015 0.67 1.075 1.35 ;
        RECT 1.1 0.54 1.16 0.73 ;
        RECT 0.195 0.67 1.485 0.73 ;
        RECT 1.425 0.6 1.485 1.35 ;
        RECT 1.51 0.54 1.57 0.66 ;
        RECT 1.425 0.6 1.57 0.66 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.8 0.06 ;
    END
  END VSS
END SDFFRHQX8

MACRO NAND4BBX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1.005 1.61 1.375 ;
        RECT 1.55 1.005 1.765 1.155 ;
        RECT 1.96 1.095 2.02 1.375 ;
        RECT 2.37 1.095 2.43 1.375 ;
        RECT 2.82 1.095 2.88 1.375 ;
        RECT 2.865 0.44 2.925 1.155 ;
        RECT 1.55 1.095 2.925 1.155 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.52 2.74 0.73 ;
        RECT 2.685 0.65 2.765 0.995 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 0.705 2.33 0.995 ;
        RECT 2.25 0.79 2.54 0.995 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.565 0.815 0.65 1.165 ;
        RECT 0.565 1.005 0.795 1.165 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.815 0.465 0.895 ;
        RECT 0.385 0.815 0.465 1.165 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.2 0.06 ;
    END
  END VSS
END NAND4BBX2

MACRO SDFFSXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSXL 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.915 1.14 1.11 ;
        RECT 1.08 0.57 1.16 0.995 ;
        RECT 1.08 0.57 1.2 0.65 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 0.57 0.54 0.63 ;
        RECT 0.46 0.57 0.52 1.22 ;
        RECT 0.46 0.57 0.54 0.73 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.425 0.645 5.485 1.025 ;
        RECT 5.32 0.965 5.485 1.025 ;
        RECT 5.615 0.585 5.675 0.705 ;
        RECT 5.835 0.625 5.965 0.705 ;
        RECT 5.425 0.645 5.97 0.705 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.585 0.815 5.945 0.895 ;
        RECT 5.865 0.805 5.945 1.025 ;
        RECT 5.755 0.815 5.945 1.025 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.98 0.585 5.06 0.98 ;
        RECT 4.98 0.585 5.165 0.705 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.635 0.625 4.765 0.705 ;
        RECT 4.685 0.625 4.765 0.96 ;
        RECT 4.685 0.88 4.88 0.96 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.815 1.965 0.895 ;
        RECT 2.105 0.29 2.165 0.875 ;
        RECT 1.715 0.815 2.165 0.875 ;
        RECT 2.105 0.29 2.77 0.35 ;
        RECT 2.71 0.29 2.77 0.47 ;
        RECT 3.09 0.35 3.15 0.47 ;
        RECT 2.71 0.41 3.15 0.47 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.2 0.06 ;
    END
  END VSS
END SDFFSXL

MACRO MX2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.495 0.42 1.63 0.48 ;
        RECT 1.525 1.05 1.585 1.48 ;
        RECT 1.57 0.42 1.63 1.11 ;
        RECT 1.57 0.98 1.74 1.11 ;
        RECT 1.525 1.05 1.995 1.11 ;
        RECT 1.935 0.39 1.995 0.53 ;
        RECT 1.57 0.47 1.995 0.53 ;
        RECT 1.935 1.05 1.995 1.48 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.815 1.315 1.105 ;
        RECT 1.18 0.95 1.315 1.105 ;
        RECT 1.235 0.815 1.47 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.63 0.54 1.13 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.34 1.29 ;
        RECT 0.64 0.91 0.7 1.29 ;
        RECT 0.26 1.23 0.7 1.29 ;
        RECT 0.64 0.91 0.76 0.97 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END MX2X4

MACRO NOR4BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BXL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.455 0.14 1.08 ;
        RECT 0.08 1.02 0.535 1.08 ;
        RECT 0.475 1.02 0.535 1.14 ;
        RECT 0.605 0.26 0.665 0.515 ;
        RECT 0.985 0.29 1.045 0.515 ;
        RECT 0.08 0.455 1.045 0.515 ;
        RECT 0.985 0.29 1.105 0.35 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.38 0.615 1.46 0.895 ;
        RECT 1.265 0.815 1.565 0.895 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 0.615 1.005 0.87 ;
        RECT 0.925 0.79 1.14 0.87 ;
        RECT 1.06 0.79 1.14 0.98 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.695 0.765 1.085 ;
        RECT 0.635 1.005 0.765 1.085 ;
        RECT 0.685 0.695 0.825 0.775 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.455 0.615 0.535 0.92 ;
        RECT 0.26 0.73 0.535 0.92 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END NOR4BXL

MACRO MXI4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X1 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.21 0.73 ;
        RECT 0.13 0.54 0.21 1.34 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.405 0.815 3.905 0.895 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.405 0.995 3.565 1.19 ;
        RECT 3.405 1.065 3.79 1.19 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.805 0.94 2.965 1.19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.585 0.805 2.705 1.085 ;
        RECT 2.405 1.005 2.705 1.085 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.59 0.815 1.765 0.895 ;
        RECT 1.685 0.815 1.765 1 ;
        RECT 1.685 0.9 1.985 1 ;
    END
  END D
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.41 0.54 0.54 ;
        RECT 0.48 0.27 0.54 0.83 ;
        RECT 0.48 0.27 1.095 0.33 ;
        RECT 1.035 0.245 1.49 0.305 ;
        RECT 1.43 0.245 1.49 0.88 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.2 0.06 ;
    END
  END VSS
END MXI4X1

MACRO OAI21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 1.14 0.705 1.48 ;
        RECT 1.06 0.79 1.14 0.92 ;
        RECT 1.06 0.86 1.3 0.92 ;
        RECT 1.195 1.14 1.255 1.48 ;
        RECT 1.24 0.6 1.3 1.2 ;
        RECT 0.645 1.14 1.3 1.2 ;
        RECT 1.325 0.54 1.385 0.66 ;
        RECT 1.24 0.6 1.385 0.66 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.96 0.54 1.3 ;
        RECT 0.46 0.96 0.7 1.04 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.345 0.78 0.94 0.86 ;
        RECT 0.86 0.78 0.94 0.92 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.4 0.76 1.48 1.2 ;
        RECT 1.4 0.79 1.54 0.92 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OAI21X2

MACRO NAND4BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX4 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.965 0.745 1.355 ;
        RECT 1.095 0.965 1.155 1.355 ;
        RECT 1.48 0.655 1.54 1.11 ;
        RECT 1.46 0.995 1.58 1.11 ;
        RECT 0.685 0.965 1.54 1.025 ;
        RECT 1.52 0.995 1.58 1.355 ;
        RECT 1.93 0.995 1.99 1.355 ;
        RECT 2.34 0.995 2.4 1.355 ;
        RECT 2.75 0.995 2.81 1.355 ;
        RECT 3.1 0.505 3.16 0.715 ;
        RECT 1.48 0.655 3.16 0.715 ;
        RECT 3.305 0.995 3.365 1.355 ;
        RECT 3.535 0.425 3.595 0.565 ;
        RECT 1.46 0.995 3.775 1.055 ;
        RECT 3.715 0.995 3.775 1.355 ;
        RECT 3.97 0.425 4.03 0.565 ;
        RECT 3.1 0.505 4.03 0.565 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.1 0.65 0.18 1.06 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 0.815 2.14 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 0.815 3.32 0.895 ;
        RECT 3.26 0.665 3.32 0.895 ;
        RECT 2.45 0.835 3.32 0.895 ;
        RECT 3.26 0.665 3.38 0.725 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.62 0.665 3.765 0.895 ;
        RECT 3.44 0.815 3.765 0.895 ;
        RECT 3.62 0.665 3.92 0.745 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.4 0.06 ;
    END
  END VSS
END NAND4BX4

MACRO TIEHI
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHI 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.9 0.14 1.4 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.6 0.06 ;
    END
  END VSS
END TIEHI

MACRO CLKINVX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX12 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.9 0.335 1.37 ;
        RECT 0.33 0.23 0.39 0.525 ;
        RECT 0.74 0.23 0.8 0.525 ;
        RECT 0.74 0.9 0.8 1.37 ;
        RECT 1.15 0.23 1.21 0.525 ;
        RECT 1.15 0.9 1.21 1.37 ;
        RECT 1.56 0.23 1.62 0.525 ;
        RECT 1.56 0.9 1.62 1.37 ;
        RECT 1.99 0.23 2.05 0.525 ;
        RECT 0.33 0.465 2.165 0.525 ;
        RECT 2.06 0.9 2.14 1.37 ;
        RECT 2.105 0.465 2.165 0.96 ;
        RECT 0.275 0.9 2.165 0.96 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.625 0.565 0.705 ;
        RECT 0.375 0.625 2.005 0.685 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END CLKINVX12

MACRO OA21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.2 0.94 1.26 1.35 ;
        RECT 1.3 0.54 1.36 0.68 ;
        RECT 1.61 0.94 1.67 1.35 ;
        RECT 1.3 0.62 1.815 0.68 ;
        RECT 1.71 0.54 1.77 0.68 ;
        RECT 1.755 0.62 1.815 1 ;
        RECT 1.755 0.79 1.94 1 ;
        RECT 1.2 0.94 1.94 1 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.63 0.14 1.13 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.63 0.605 0.71 ;
        RECT 0.435 0.63 0.605 0.895 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.72 0.61 0.8 0.87 ;
        RECT 0.72 0.79 0.94 0.87 ;
        RECT 0.86 0.79 0.94 0.97 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END OA21X4

MACRO AOI221XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221XL 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.965 0.475 1.025 0.7 ;
        RECT 1.715 0.475 1.775 0.7 ;
        RECT 0.965 0.64 1.88 0.7 ;
        RECT 1.82 0.64 1.88 1.21 ;
        RECT 1.82 0.79 1.94 0.92 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.69 0.815 0.965 0.955 ;
        RECT 0.69 0.875 1.13 0.955 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 0.815 1.325 1.085 ;
        RECT 1.23 0.815 1.54 0.895 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.835 0.395 1.085 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 0.8 1.72 1.085 ;
        RECT 1.425 1.005 1.72 1.085 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.245 0.565 0.325 ;
        RECT 0.47 0.245 0.565 0.735 ;
        RECT 0.47 0.655 0.59 0.735 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2 0.06 ;
    END
  END VSS
END AOI221XL

MACRO DLY2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY2X1 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.415 0.14 1.175 ;
        RECT 0.08 1.115 0.33 1.175 ;
        RECT 0.27 0.355 0.33 0.475 ;
        RECT 0.08 0.415 0.33 0.475 ;
        RECT 0.27 1.115 0.33 1.395 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.625 1.52 1.08 ;
        RECT 1.46 0.6 1.54 0.73 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.4 0.06 ;
    END
  END VSS
END DLY2X1

MACRO OAI31X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X4 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.915 1.125 0.975 1.405 ;
        RECT 2.165 1.125 2.225 1.405 ;
        RECT 0.915 1.125 3.135 1.185 ;
        RECT 3.06 0.485 3.12 1.185 ;
        RECT 3.075 0.98 3.135 1.405 ;
        RECT 3.06 0.98 3.14 1.11 ;
        RECT 3.06 0.485 3.265 0.595 ;
        RECT 3.06 1.05 3.545 1.11 ;
        RECT 3.485 1.015 3.545 1.405 ;
        RECT 3.06 0.535 3.6 0.595 ;
        RECT 3.54 0.485 3.675 0.545 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.22 0.8 3.705 0.88 ;
        RECT 3.425 0.8 3.705 0.895 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.815 0.365 0.935 ;
        RECT 0.235 0.875 0.665 0.935 ;
        RECT 0.605 0.875 0.665 1.025 ;
        RECT 1.425 0.885 1.545 1.025 ;
        RECT 2.76 0.855 2.82 1.025 ;
        RECT 0.605 0.965 2.82 1.025 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 0.655 0.825 0.715 ;
        RECT 0.765 0.655 0.825 0.865 ;
        RECT 1.265 0.725 1.325 0.865 ;
        RECT 0.765 0.805 1.325 0.865 ;
        RECT 1.265 0.725 1.705 0.785 ;
        RECT 1.645 0.725 1.705 0.865 ;
        RECT 2.26 0.6 2.32 0.865 ;
        RECT 1.645 0.805 2.32 0.865 ;
        RECT 2.26 0.6 2.34 0.745 ;
        RECT 2.26 0.625 2.565 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.625 1.165 0.705 ;
        RECT 0.925 0.645 1.165 0.705 ;
        RECT 1.105 0.565 1.865 0.625 ;
        RECT 1.805 0.565 1.865 0.705 ;
        RECT 1.805 0.645 2.115 0.705 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4 0.06 ;
    END
  END VSS
END OAI31X4

MACRO TLATNTSCAX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX12 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.235 0.35 4.295 0.66 ;
        RECT 4.235 0.87 4.295 1.42 ;
        RECT 4.235 0.87 4.3 0.925 ;
        RECT 4.26 0.605 4.32 0.92 ;
        RECT 4.26 0.79 4.34 0.92 ;
        RECT 4.645 0.35 4.705 1.42 ;
        RECT 5.055 0.35 5.115 1.42 ;
        RECT 5.465 0.35 5.525 1.42 ;
        RECT 5.83 0.79 5.89 1.01 ;
        RECT 5.875 0.35 5.935 0.85 ;
        RECT 4.26 0.79 5.935 0.85 ;
        RECT 5.875 0.95 5.935 1.42 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.745 0.73 ;
        RECT 0.665 0.45 0.745 0.945 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.45 0.54 0.945 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.060 0.48 0.14 0.895 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END TLATNTSCAX12

MACRO NAND3BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BXL 0 0 ;
  SIZE 1.00 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 1.005 0.14 1.085 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.725 0.765 0.81 0.895 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.33 0.41 0.41 0.515 ;
        RECT 0.33 0.46 0.465 0.515 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.18 0.6 0.27 0.705 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.00 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.00 0.06 ;
    END
  END VSS
END NAND3BXL

MACRO EDFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFX4 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.245 1.05 5.305 1.44 ;
        RECT 5.26 0.57 5.32 1.11 ;
        RECT 5.26 0.98 5.34 1.11 ;
        RECT 5.245 1.05 5.715 1.11 ;
        RECT 5.1 0.57 5.69 0.63 ;
        RECT 5.655 1.05 5.715 1.44 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.425 1.05 4.485 1.44 ;
        RECT 4.46 0.57 4.52 1.11 ;
        RECT 4.46 0.98 4.54 1.11 ;
        RECT 4.16 0.57 4.75 0.63 ;
        RECT 4.425 1.05 4.895 1.11 ;
        RECT 4.835 1.05 4.895 1.44 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.645 0.815 4.145 0.895 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.885 0.815 3.165 0.895 ;
        RECT 3.045 0.815 3.165 1.115 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.765 0.34 1.265 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.4 0.06 ;
    END
  END VSS
END EDFFX4

MACRO OAI222X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.695 1.19 0.755 1.47 ;
        RECT 1.44 0.37 1.5 0.51 ;
        RECT 1.495 1.19 1.555 1.47 ;
        RECT 1.44 0.45 1.72 0.51 ;
        RECT 1.66 0.45 1.72 1.25 ;
        RECT 1.66 0.98 1.74 1.25 ;
        RECT 0.695 1.19 1.74 1.25 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 0.68 0.83 1.09 ;
        RECT 0.66 0.79 0.83 1.09 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.68 0.34 1.18 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.59 1.34 1.09 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 0.68 0.52 1.06 ;
        RECT 0.46 0.98 0.54 1.16 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.48 0.61 1.56 1.09 ;
        RECT 1.46 0.79 1.56 1.09 ;
    END
  END C1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.45 1.14 0.95 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OAI222X1

MACRO SDFFRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX2 0 0 ;
  SIZE 5.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 0.42 0.335 1.005 ;
        RECT 0.26 0.925 0.34 1.315 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.78 0.645 4.84 0.915 ;
        RECT 5.035 0.625 5.165 0.705 ;
        RECT 4.78 0.645 5.2 0.705 ;
        RECT 5.14 0.655 5.475 0.715 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.195 0.815 5.61 0.925 ;
        RECT 5.14 0.845 5.61 0.925 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.6 4.34 0.73 ;
        RECT 4.26 0.6 4.52 0.68 ;
        RECT 4.44 0.6 4.52 0.87 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.48 0.79 1.665 0.995 ;
        RECT 1.48 0.815 1.855 0.995 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 0.66 0.74 0.92 ;
        RECT 0.66 0.66 0.74 1.095 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.8 0.06 ;
    END
  END VSS
END SDFFRHQX2

MACRO CLKMX2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.495 0.42 1.63 0.48 ;
        RECT 1.525 1.05 1.585 1.48 ;
        RECT 1.57 0.42 1.63 1.11 ;
        RECT 1.57 0.98 1.74 1.11 ;
        RECT 1.525 1.05 1.995 1.11 ;
        RECT 1.935 0.39 1.995 0.53 ;
        RECT 1.57 0.47 1.995 0.53 ;
        RECT 1.935 1.05 1.995 1.48 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.815 1.315 1.105 ;
        RECT 1.18 0.95 1.315 1.105 ;
        RECT 1.235 0.815 1.47 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.63 0.54 1.13 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.34 1.29 ;
        RECT 0.64 0.91 0.7 1.29 ;
        RECT 0.26 1.23 0.7 1.29 ;
        RECT 0.64 0.91 0.76 0.97 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END CLKMX2X4

MACRO EDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRX2 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.065 0.54 7.145 1.11 ;
        RECT 7.06 0.98 7.145 1.11 ;
        RECT 7.06 1.03 7.215 1.11 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.675 0.54 6.755 1.14 ;
        RECT 6.625 1.06 6.755 1.14 ;
        RECT 6.675 0.79 6.94 0.92 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.285 0.635 6.365 1.085 ;
        RECT 6.235 1.005 6.365 1.085 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.75 2.74 1.25 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.005 0.765 1.085 ;
        RECT 0.705 0.73 0.765 1.15 ;
        RECT 1.305 0.77 1.365 1.15 ;
        RECT 0.705 1.09 1.365 1.15 ;
        RECT 1.305 0.77 1.48 0.83 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.88 ;
        RECT 0.26 0.6 0.56 0.73 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 7.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 7.8 0.06 ;
    END
  END VSS
END EDFFTRX2

MACRO CLKAND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X6 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 0.275 1.855 0.585 ;
        RECT 1.85 0.86 1.91 1.37 ;
        RECT 2.205 0.275 2.265 0.585 ;
        RECT 2.26 0.86 2.32 1.37 ;
        RECT 2.46 0.525 2.52 0.92 ;
        RECT 2.46 0.79 2.54 0.92 ;
        RECT 1.85 0.86 2.73 0.92 ;
        RECT 2.615 0.275 2.675 0.585 ;
        RECT 1.795 0.525 2.675 0.585 ;
        RECT 2.67 0.86 2.73 1.37 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.54 0.785 0.66 0.895 ;
        RECT 1.07 0.785 1.19 0.895 ;
        RECT 0.54 0.815 1.19 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 0.645 0.365 0.705 ;
        RECT 0.235 0.625 1.535 0.685 ;
        RECT 1.475 0.625 1.535 0.745 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.8 0.06 ;
    END
  END VSS
END CLKAND2X6

MACRO OA21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.2 0.67 1.26 1.455 ;
        RECT 1.26 0.6 1.34 0.73 ;
        RECT 1.28 0.57 1.495 0.63 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.56 0.34 1.06 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.785 0.54 0.925 ;
        RECT 0.625 0.59 0.705 0.865 ;
        RECT 0.46 0.785 0.705 0.865 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.22 0.94 0.72 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END OA21X2

MACRO OAI31X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X2 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.91 1.185 0.97 1.305 ;
        RECT 1.46 0.98 1.54 1.245 ;
        RECT 1.46 1.05 1.715 1.245 ;
        RECT 0.91 1.185 1.715 1.245 ;
        RECT 1.655 1.05 1.715 1.435 ;
        RECT 1.7 0.545 1.76 1.11 ;
        RECT 1.7 0.545 1.875 0.605 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.945 0.915 1.165 1.085 ;
        RECT 0.89 1.005 1.165 1.085 ;
        RECT 0.945 0.915 1.3 0.995 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.755 0.74 0.92 ;
        RECT 0.495 0.755 1.235 0.815 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.335 0.595 0.395 0.795 ;
        RECT 0.335 0.595 1.46 0.655 ;
        RECT 1.4 0.6 1.54 0.82 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.705 1.94 1.205 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.2 0.06 ;
    END
  END VSS
END OAI31X2

MACRO EDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX1 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.1 0.535 3.18 1.09 ;
        RECT 3.06 0.79 3.18 1.09 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.835 0.305 3.895 0.905 ;
        RECT 4.185 0.625 4.245 0.745 ;
        RECT 3.835 0.305 4.36 0.365 ;
        RECT 4.3 0.305 4.36 0.685 ;
        RECT 4.185 0.625 4.765 0.685 ;
        RECT 4.555 0.625 4.765 0.715 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.375 0.785 4.455 0.97 ;
        RECT 4.375 0.815 4.77 0.935 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.73 0.34 1.23 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5 0.06 ;
    END
  END VSS
END EDFFHQX1

MACRO SDFFSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX2 0 0 ;
  SIZE 9.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.46 0.6 8.54 0.73 ;
        RECT 8.46 0.67 8.7 0.73 ;
        RECT 8.64 0.57 8.7 1.305 ;
        RECT 8.64 0.57 8.76 0.63 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.06 0.98 8.2 1.11 ;
        RECT 8.12 0.54 8.2 1.305 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.635 0.73 7.715 1.085 ;
        RECT 7.635 0.95 7.86 1.085 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 0.625 3.365 0.8 ;
        RECT 3.205 0.675 3.61 0.755 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.525 1.74 1.025 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.28 0.6 1.36 0.87 ;
        RECT 1.28 0.6 1.54 0.68 ;
        RECT 1.46 0.6 1.54 0.73 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.715 0.685 0.92 ;
        RECT 0.605 0.715 0.685 1.07 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.655 0.23 0.715 0.615 ;
        RECT 0.28 0.555 0.775 0.615 ;
        RECT 0.74 0.56 0.86 0.62 ;
        RECT 0.655 0.23 1.18 0.29 ;
        RECT 1.12 0.23 1.18 1.03 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 9.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 9.4 0.06 ;
    END
  END VSS
END SDFFSRX2

MACRO OA22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 1.05 1.3 1.44 ;
        RECT 1.49 0.44 1.61 0.5 ;
        RECT 1.65 1.05 1.71 1.44 ;
        RECT 1.56 0.46 2.005 0.52 ;
        RECT 1.945 0.41 2.005 1.11 ;
        RECT 1.945 0.98 2.14 1.11 ;
        RECT 1.24 1.05 2.14 1.11 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.78 1.08 1.06 ;
        RECT 1.06 0.98 1.14 1.22 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 0.72 0.56 1.2 ;
        RECT 0.46 0.88 0.56 1.2 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.72 0.34 1.22 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.72 0.74 1.22 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 2.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 2.4 0.06 ;
    END
  END VSS
END OA22X4

MACRO CLKAND2X3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X3 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.065 0.445 1.185 0.505 ;
        RECT 1.155 0.945 1.215 1.335 ;
        RECT 1.46 0.495 1.54 1.005 ;
        RECT 1.155 0.945 1.625 1.005 ;
        RECT 1.505 0.415 1.565 0.555 ;
        RECT 1.125 0.495 1.565 0.555 ;
        RECT 1.565 0.945 1.625 1.335 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.805 0.57 0.925 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.215 0.625 0.805 0.705 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.8 0.06 ;
    END
  END VSS
END CLKAND2X3

MACRO EDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFX2 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.66 0.6 4.74 0.73 ;
        RECT 4.68 0.505 4.74 1.355 ;
        RECT 4.68 0.505 4.815 0.565 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.225 0.505 4.345 0.565 ;
        RECT 4.235 0.505 4.295 1.355 ;
        RECT 4.235 0.505 4.345 0.705 ;
        RECT 4.235 0.625 4.365 0.705 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.805 1.25 2.865 1.485 ;
        RECT 2.745 1.425 2.865 1.485 ;
        RECT 2.955 0.665 3.075 0.725 ;
        RECT 3.015 0.665 3.075 1.31 ;
        RECT 3.86 0.775 3.92 1.31 ;
        RECT 2.805 1.25 3.92 1.31 ;
        RECT 3.835 0.775 3.955 0.895 ;
        RECT 3.835 0.815 3.965 0.895 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.395 0.64 3.54 0.725 ;
        RECT 3.46 0.64 3.54 1.04 ;
        RECT 3.395 0.64 3.575 0.72 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.775 0.315 1.025 ;
        RECT 0.325 0.62 0.405 0.895 ;
        RECT 0.23 0.775 0.405 0.895 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END EDFFX2

MACRO DLY3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY3X1 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.635 0.54 2.695 0.895 ;
        RECT 2.635 0.815 2.89 0.895 ;
        RECT 2.83 0.815 2.89 1.29 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 0.76 1.935 1.065 ;
        RECT 1.66 0.79 1.935 1.065 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.8 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.8 0.06 ;
    END
  END VSS
END DLY3X1

MACRO OAI222X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.155 0.835 1.275 ;
        RECT 1.445 1.155 1.505 1.275 ;
        RECT 2.365 1.155 2.425 1.275 ;
        RECT 3.22 1.155 3.28 1.275 ;
        RECT 3.835 0.535 3.895 0.675 ;
        RECT 4.005 1.155 4.065 1.275 ;
        RECT 4.245 0.535 4.305 0.675 ;
        RECT 4.63 1.155 4.69 1.275 ;
        RECT 4.655 0.535 4.715 0.675 ;
        RECT 3.835 0.615 5.125 0.675 ;
        RECT 5.06 0.615 5.12 1.215 ;
        RECT 0.775 1.155 5.12 1.215 ;
        RECT 5.065 0.535 5.125 0.92 ;
        RECT 5.06 0.79 5.14 0.92 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 0.935 0.365 1.055 ;
        RECT 1.065 0.935 1.185 1.055 ;
        RECT 1.66 0.79 1.74 1.055 ;
        RECT 0.305 0.995 1.74 1.055 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.73 0.835 3.94 0.895 ;
        RECT 3.86 0.79 3.94 1.055 ;
        RECT 4.35 0.935 4.47 1.055 ;
        RECT 4.865 0.895 4.925 1.055 ;
        RECT 3.86 0.995 4.925 1.055 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.085 0.895 2.145 1.055 ;
        RECT 2.685 0.935 2.805 1.055 ;
        RECT 3.46 0.79 3.52 1.055 ;
        RECT 2.085 0.995 3.52 1.055 ;
        RECT 3.46 0.79 3.54 0.92 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 0.775 0.965 0.895 ;
        RECT 0.67 0.775 1.47 0.835 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.04 0.775 4.765 0.835 ;
        RECT 4.635 0.775 4.765 0.895 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.435 0.775 2.585 0.895 ;
        RECT 2.435 0.775 3.18 0.835 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END OAI222X4

MACRO INVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.465 0.54 0.535 0.71 ;
#        RECT 0.46 0.72 0.54 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.6 0.175 0.8 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 0.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 0.6 0.06 ;
    END
  END VSS
END INVX2

MACRO TLATNSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRXL 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.545 0.94 1.11 ;
        RECT 0.86 1.03 1.055 1.11 ;
        RECT 0.975 0.505 1.055 0.625 ;
        RECT 0.86 0.545 1.055 0.625 ;
        RECT 0.975 1.03 1.055 1.175 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.325 0.73 ;
        RECT 0.245 0.54 0.325 1.02 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.83 4.34 1.26 ;
        RECT 4.26 0.83 4.41 1.11 ;
    END
  END GN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 0.345 3.79 0.405 ;
        RECT 3.73 0.345 3.79 0.92 ;
        RECT 3.66 0.79 3.79 0.92 ;
        RECT 3.66 0.86 4.16 0.92 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 0.665 3.025 1.01 ;
        RECT 2.945 0.665 3.18 0.92 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.285 0.885 1.365 1.275 ;
        RECT 1.175 1.195 1.365 1.275 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 4.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 4.6 0.06 ;
    END
  END VSS
END TLATNSRXL

MACRO MXI2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 0.73 ;
        RECT 0.28 0.48 0.34 1.265 ;
        RECT 0.28 0.48 0.52 0.54 ;
        RECT 0.28 1.205 0.605 1.265 ;
        RECT 0.545 1.205 0.605 1.325 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 0.8 1.14 0.88 ;
        RECT 1.06 0.8 1.14 1.11 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.77 0.98 0.96 1.2 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.74 0.14 0.92 ;
        RECT 0.1 0.84 0.18 1.2 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.4 0.06 ;
    END
  END VSS
END MXI2XL

MACRO NAND4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.41 1.14 0.635 ;
        RECT 1.08 0.41 1.14 1.015 ;
        RECT 0.365 0.955 1.14 1.015 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.355 0.34 0.855 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.355 0.54 0.855 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.355 0.74 0.855 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.355 0.94 0.855 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 1.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 1.2 0.06 ;
    END
  END VSS
END NAND4XL

MACRO DFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX8 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.04 0.67 5.19 0.94 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.63 0.67 4.71 0.92 ;
        RECT 4.63 0.785 4.94 0.92 ;
        RECT 4.86 0.785 4.94 0.94 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 0.73 ;
        RECT 0.08 0.54 0.14 1.345 ;
        RECT 0.06 0.67 0.55 0.73 ;
        RECT 0.49 0.54 0.55 1.345 ;
        RECT 0.9 0.54 0.96 1.345 ;
        RECT 0.49 0.6 1.37 0.66 ;
        RECT 1.31 0.54 1.37 1.345 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 5.4 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 5.4 0.06 ;
    END
  END VSS
END DFFHQX8

MACRO EDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX4 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.02 0.57 3.14 0.63 ;
        RECT 3.08 0.57 3.14 1.085 ;
        RECT 3.035 1.005 3.225 1.085 ;
        RECT 3.165 1.005 3.225 1.16 ;
        RECT 3.17 1.125 3.725 1.185 ;
        RECT 3.78 0.57 3.84 0.81 ;
        RECT 3.08 0.75 3.84 0.81 ;
        RECT 3.78 0.57 3.9 0.63 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.92 0.245 4.98 0.915 ;
        RECT 4.92 0.245 5.36 0.305 ;
        RECT 5.3 0.245 5.36 0.685 ;
        RECT 5.24 0.625 5.36 0.685 ;
        RECT 5.3 0.485 5.895 0.545 ;
        RECT 5.835 0.485 5.895 0.705 ;
        RECT 5.835 0.625 5.965 0.705 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.655 0.645 5.735 0.95 ;
        RECT 5.46 0.79 5.735 0.95 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.81 0.34 1.31 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 6.2 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 6.2 0.06 ;
    END
  END VSS
END EDFFHQX4

MACRO TLATNCAX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX4 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.9 0.7 1.02 ;
        RECT 0.66 0.51 0.72 0.96 ;
        RECT 0.66 0.79 0.74 0.96 ;
        RECT 0.66 0.57 1.105 0.63 ;
        RECT 0.64 0.9 1.14 0.96 ;
        RECT 1.055 0.55 1.175 0.61 ;
        RECT 1.08 0.93 1.2 0.99 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.95 0.78 3.03 1.06 ;
        RECT 2.95 0.78 3.25 0.895 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.33 0.65 0.41 0.97 ;
        RECT 0.46 0.6 0.54 0.73 ;
        RECT 0.33 0.65 0.54 0.73 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 1.65 3.6 1.71 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 0.00 3.6 0.06 ;
    END
  END VSS
END TLATNCAX4

MACRO MEM1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM1 0 0 ;
  SIZE 426.965 BY 114.215 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.000 77.64 12.660 78.3 ;
      LAYER Metal6 ;
        RECT 12.000 77.64 12.660 78.3 ;
      LAYER Metal3 ;
        RECT 12.000 77.64 12.660 78.3 ;
      LAYER Metal4 ;
        RECT 12.000 77.64 12.660 78.3 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.000 71.52 12.660 72.18 ;
      LAYER Metal6 ;
        RECT 12.000 71.52 12.660 72.18 ;
      LAYER Metal3 ;
        RECT 12.000 71.52 12.660 72.18 ;
      LAYER Metal4 ;
        RECT 12.000 71.52 12.660 72.18 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.000 68.42 12.660 69.08 ;
      LAYER Metal6 ;
        RECT 12.000 68.42 12.660 69.08 ;
      LAYER Metal3 ;
        RECT 12.000 68.42 12.660 69.08 ;
      LAYER Metal4 ;
        RECT 12.000 68.42 12.660 69.08 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.000 62.3 12.660 62.96 ;
      LAYER Metal6 ;
        RECT 12.000 62.3 12.660 62.96 ;
      LAYER Metal3 ;
        RECT 12.000 62.3 12.660 62.96 ;
      LAYER Metal4 ;
        RECT 12.000 62.3 12.660 62.96 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.000 59.28 12.660 59.94 ;
      LAYER Metal6 ;
        RECT 12.000 59.28 12.660 59.94 ;
      LAYER Metal3 ;
        RECT 12.000 59.28 12.660 59.94 ;
      LAYER Metal4 ;
        RECT 12.000 59.28 12.660 59.94 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.000 56.18 12.660 56.84 ;
      LAYER Metal6 ;
        RECT 12.000 56.18 12.660 56.84 ;
      LAYER Metal3 ;
        RECT 12.000 56.18 12.660 56.84 ;
      LAYER Metal4 ;
        RECT 12.000 56.18 12.660 56.84 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.000 50.06 12.660 50.72 ;
      LAYER Metal6 ;
        RECT 12.000 50.06 12.660 50.72 ;
      LAYER Metal3 ;
        RECT 12.000 50.06 12.660 50.72 ;
      LAYER Metal4 ;
        RECT 12.000 50.06 12.660 50.72 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.000 47.04 12.660 47.7 ;
      LAYER Metal6 ;
        RECT 12.000 47.04 12.660 47.7 ;
      LAYER Metal3 ;
        RECT 12.000 47.04 12.660 47.7 ;
      LAYER Metal4 ;
        RECT 12.000 47.04 12.660 47.7 ;
    END
  END A[7]
  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 228.435 12 229.095 12.66 ;
      LAYER Metal6 ;
        RECT 228.435 12 229.095 12.66 ;
      LAYER Metal3 ;
        RECT 228.435 12 229.095 12.66 ;
      LAYER Metal4 ;
        RECT 228.435 12 229.095 12.66 ;
    END
  END CE
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal5 ;
        RECT 238.18 12 238.84 12.66 ;
      LAYER Metal6 ;
        RECT 238.18 12 238.84 12.66 ;
      LAYER Metal3 ;
        RECT 238.18 12 238.84 12.66 ;
      LAYER Metal4 ;
        RECT 238.18 12 238.84 12.66 ;
    END
  END CK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 20.48 12 21.14 12.66 ;
      LAYER Metal6 ;
        RECT 20.48 12 21.14 12.66 ;
      LAYER Metal3 ;
        RECT 20.48 12 21.14 12.66 ;
      LAYER Metal4 ;
        RECT 20.48 12 21.14 12.66 ;
    END
  END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 129 12 129.66 12.66 ;
      LAYER Metal6 ;
        RECT 129 12 129.66 12.66 ;
      LAYER Metal3 ;
        RECT 129 12 129.66 12.66 ;
      LAYER Metal4 ;
        RECT 129 12 129.66 12.66 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 137.04 12 137.7 12.66 ;
      LAYER Metal6 ;
        RECT 137.04 12 137.7 12.66 ;
      LAYER Metal3 ;
        RECT 137.04 12 137.7 12.66 ;
      LAYER Metal4 ;
        RECT 137.04 12 137.7 12.66 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 151.34 12 152 12.66 ;
      LAYER Metal6 ;
        RECT 151.34 12 152 12.66 ;
      LAYER Metal3 ;
        RECT 151.34 12 152 12.66 ;
      LAYER Metal4 ;
        RECT 151.34 12 152 12.66 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 159.38 12 160.04 12.66 ;
      LAYER Metal6 ;
        RECT 159.38 12 160.04 12.66 ;
      LAYER Metal3 ;
        RECT 159.38 12 160.04 12.66 ;
      LAYER Metal4 ;
        RECT 159.38 12 160.04 12.66 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 172.62 12 173.28 12.66 ;
      LAYER Metal6 ;
        RECT 172.62 12 173.28 12.66 ;
      LAYER Metal3 ;
        RECT 172.62 12 173.28 12.66 ;
      LAYER Metal4 ;
        RECT 172.62 12 173.28 12.66 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 180.66 12 181.32 12.66 ;
      LAYER Metal6 ;
        RECT 180.66 12 181.32 12.66 ;
      LAYER Metal3 ;
        RECT 180.66 12 181.32 12.66 ;
      LAYER Metal4 ;
        RECT 180.66 12 181.32 12.66 ;
    END
  END D[15]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 245.645 12 246.305 12.66 ;
      LAYER Metal6 ;
        RECT 245.645 12 246.305 12.66 ;
      LAYER Metal3 ;
        RECT 245.645 12 246.305 12.66 ;
      LAYER Metal4 ;
        RECT 245.645 12 246.305 12.66 ;
    END
  END D[16]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 253.685 12 254.345 12.66 ;
      LAYER Metal6 ;
        RECT 253.685 12 254.345 12.66 ;
      LAYER Metal3 ;
        RECT 253.685 12 254.345 12.66 ;
      LAYER Metal4 ;
        RECT 253.685 12 254.345 12.66 ;
    END
  END D[17]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 266.925 12 267.585 12.66 ;
      LAYER Metal6 ;
        RECT 266.925 12 267.585 12.66 ;
      LAYER Metal3 ;
        RECT 266.925 12 267.585 12.66 ;
      LAYER Metal4 ;
        RECT 266.925 12 267.585 12.66 ;
    END
  END D[18]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 274.965 12 275.625 12.66 ;
      LAYER Metal6 ;
        RECT 274.965 12 275.625 12.66 ;
      LAYER Metal3 ;
        RECT 274.965 12 275.625 12.66 ;
      LAYER Metal4 ;
        RECT 274.965 12 275.625 12.66 ;
    END
  END D[19]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 28.52 12 29.18 12.66 ;
      LAYER Metal6 ;
        RECT 28.52 12 29.18 12.66 ;
      LAYER Metal3 ;
        RECT 28.52 12 29.18 12.66 ;
      LAYER Metal4 ;
        RECT 28.52 12 29.18 12.66 ;
    END
  END D[1]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 289.265 12 289.925 12.66 ;
      LAYER Metal6 ;
        RECT 289.265 12 289.925 12.66 ;
      LAYER Metal3 ;
        RECT 289.265 12 289.925 12.66 ;
      LAYER Metal4 ;
        RECT 289.265 12 289.925 12.66 ;
    END
  END D[20]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 297.305 12 297.965 12.66 ;
      LAYER Metal6 ;
        RECT 297.305 12 297.965 12.66 ;
      LAYER Metal3 ;
        RECT 297.305 12 297.965 12.66 ;
      LAYER Metal4 ;
        RECT 297.305 12 297.965 12.66 ;
    END
  END D[21]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 310.545 12 311.205 12.66 ;
      LAYER Metal6 ;
        RECT 310.545 12 311.205 12.66 ;
      LAYER Metal3 ;
        RECT 310.545 12 311.205 12.66 ;
      LAYER Metal4 ;
        RECT 310.545 12 311.205 12.66 ;
    END
  END D[22]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 318.585 12 319.245 12.66 ;
      LAYER Metal6 ;
        RECT 318.585 12 319.245 12.66 ;
      LAYER Metal3 ;
        RECT 318.585 12 319.245 12.66 ;
      LAYER Metal4 ;
        RECT 318.585 12 319.245 12.66 ;
    END
  END D[23]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 332.885 12 333.545 12.66 ;
      LAYER Metal6 ;
        RECT 332.885 12 333.545 12.66 ;
      LAYER Metal3 ;
        RECT 332.885 12 333.545 12.66 ;
      LAYER Metal4 ;
        RECT 332.885 12 333.545 12.66 ;
    END
  END D[24]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 340.925 12 341.585 12.66 ;
      LAYER Metal6 ;
        RECT 340.925 12 341.585 12.66 ;
      LAYER Metal3 ;
        RECT 340.925 12 341.585 12.66 ;
      LAYER Metal4 ;
        RECT 340.925 12 341.585 12.66 ;
    END
  END D[25]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 354.165 12 354.825 12.66 ;
      LAYER Metal6 ;
        RECT 354.165 12 354.825 12.66 ;
      LAYER Metal3 ;
        RECT 354.165 12 354.825 12.66 ;
      LAYER Metal4 ;
        RECT 354.165 12 354.825 12.66 ;
    END
  END D[26]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 362.205 12 362.865 12.66 ;
      LAYER Metal6 ;
        RECT 362.205 12 362.865 12.66 ;
      LAYER Metal3 ;
        RECT 362.205 12 362.865 12.66 ;
      LAYER Metal4 ;
        RECT 362.205 12 362.865 12.66 ;
    END
  END D[27]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.505 12 377.165 12.66 ;
      LAYER Metal6 ;
        RECT 376.505 12 377.165 12.66 ;
      LAYER Metal3 ;
        RECT 376.505 12 377.165 12.66 ;
      LAYER Metal4 ;
        RECT 376.505 12 377.165 12.66 ;
    END
  END D[28]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.545 12 385.205 12.66 ;
      LAYER Metal6 ;
        RECT 384.545 12 385.205 12.66 ;
      LAYER Metal3 ;
        RECT 384.545 12 385.205 12.66 ;
      LAYER Metal4 ;
        RECT 384.545 12 385.205 12.66 ;
    END
  END D[29]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 41.76 12 42.42 12.66 ;
      LAYER Metal6 ;
        RECT 41.76 12 42.42 12.66 ;
      LAYER Metal3 ;
        RECT 41.76 12 42.42 12.66 ;
      LAYER Metal4 ;
        RECT 41.76 12 42.42 12.66 ;
    END
  END D[2]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 397.785 12 398.445 12.66 ;
      LAYER Metal6 ;
        RECT 397.785 12 398.445 12.66 ;
      LAYER Metal3 ;
        RECT 397.785 12 398.445 12.66 ;
      LAYER Metal4 ;
        RECT 397.785 12 398.445 12.66 ;
    END
  END D[30]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 405.825 12 406.485 12.66 ;
      LAYER Metal6 ;
        RECT 405.825 12 406.485 12.66 ;
      LAYER Metal3 ;
        RECT 405.825 12 406.485 12.66 ;
      LAYER Metal4 ;
        RECT 405.825 12 406.485 12.66 ;
    END
  END D[31]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 49.8 12 50.46 12.66 ;
      LAYER Metal6 ;
        RECT 49.8 12 50.46 12.66 ;
      LAYER Metal3 ;
        RECT 49.8 12 50.46 12.66 ;
      LAYER Metal4 ;
        RECT 49.8 12 50.46 12.66 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.1 12 64.76 12.66 ;
      LAYER Metal6 ;
        RECT 64.1 12 64.76 12.66 ;
      LAYER Metal3 ;
        RECT 64.1 12 64.76 12.66 ;
      LAYER Metal4 ;
        RECT 64.1 12 64.76 12.66 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.14 12 72.8 12.66 ;
      LAYER Metal6 ;
        RECT 72.14 12 72.8 12.66 ;
      LAYER Metal3 ;
        RECT 72.14 12 72.8 12.66 ;
      LAYER Metal4 ;
        RECT 72.14 12 72.8 12.66 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.38 12 86.04 12.66 ;
      LAYER Metal6 ;
        RECT 85.38 12 86.04 12.66 ;
      LAYER Metal3 ;
        RECT 85.38 12 86.04 12.66 ;
      LAYER Metal4 ;
        RECT 85.38 12 86.04 12.66 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.42 12 94.08 12.66 ;
      LAYER Metal6 ;
        RECT 93.42 12 94.08 12.66 ;
      LAYER Metal3 ;
        RECT 93.42 12 94.08 12.66 ;
      LAYER Metal4 ;
        RECT 93.42 12 94.08 12.66 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.72 12 108.38 12.66 ;
      LAYER Metal6 ;
        RECT 107.72 12 108.38 12.66 ;
      LAYER Metal3 ;
        RECT 107.72 12 108.38 12.66 ;
      LAYER Metal4 ;
        RECT 107.72 12 108.38 12.66 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 115.76 12 116.42 12.66 ;
      LAYER Metal6 ;
        RECT 115.76 12 116.42 12.66 ;
      LAYER Metal3 ;
        RECT 115.76 12 116.42 12.66 ;
      LAYER Metal4 ;
        RECT 115.76 12 116.42 12.66 ;
    END
  END D[9]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 23.06 12 23.72 12.66 ;
      LAYER Metal6 ;
        RECT 23.06 12 23.72 12.66 ;
      LAYER Metal3 ;
        RECT 23.06 12 23.72 12.66 ;
      LAYER Metal4 ;
        RECT 23.06 12 23.72 12.66 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.58 12 132.24 12.66 ;
      LAYER Metal6 ;
        RECT 131.58 12 132.24 12.66 ;
      LAYER Metal3 ;
        RECT 131.58 12 132.24 12.66 ;
      LAYER Metal4 ;
        RECT 131.58 12 132.24 12.66 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 134.46 12 135.12 12.66 ;
      LAYER Metal6 ;
        RECT 134.46 12 135.12 12.66 ;
      LAYER Metal3 ;
        RECT 134.46 12 135.12 12.66 ;
      LAYER Metal4 ;
        RECT 134.46 12 135.12 12.66 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.92 12 154.58 12.66 ;
      LAYER Metal6 ;
        RECT 153.92 12 154.58 12.66 ;
      LAYER Metal3 ;
        RECT 153.92 12 154.58 12.66 ;
      LAYER Metal4 ;
        RECT 153.92 12 154.58 12.66 ;
    END
  END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 156.8 12 157.46 12.66 ;
      LAYER Metal6 ;
        RECT 156.8 12 157.46 12.66 ;
      LAYER Metal3 ;
        RECT 156.8 12 157.46 12.66 ;
      LAYER Metal4 ;
        RECT 156.8 12 157.46 12.66 ;
    END
  END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.2 12 175.86 12.66 ;
      LAYER Metal6 ;
        RECT 175.2 12 175.86 12.66 ;
      LAYER Metal3 ;
        RECT 175.2 12 175.86 12.66 ;
      LAYER Metal4 ;
        RECT 175.2 12 175.86 12.66 ;
    END
  END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.08 12 178.74 12.66 ;
      LAYER Metal6 ;
        RECT 178.08 12 178.74 12.66 ;
      LAYER Metal3 ;
        RECT 178.08 12 178.74 12.66 ;
      LAYER Metal4 ;
        RECT 178.08 12 178.74 12.66 ;
    END
  END Q[15]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 248.225 12 248.885 12.66 ;
      LAYER Metal6 ;
        RECT 248.225 12 248.885 12.66 ;
      LAYER Metal3 ;
        RECT 248.225 12 248.885 12.66 ;
      LAYER Metal4 ;
        RECT 248.225 12 248.885 12.66 ;
    END
  END Q[16]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 251.105 12 251.765 12.66 ;
      LAYER Metal6 ;
        RECT 251.105 12 251.765 12.66 ;
      LAYER Metal3 ;
        RECT 251.105 12 251.765 12.66 ;
      LAYER Metal4 ;
        RECT 251.105 12 251.765 12.66 ;
    END
  END Q[17]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 269.505 12 270.165 12.66 ;
      LAYER Metal6 ;
        RECT 269.505 12 270.165 12.66 ;
      LAYER Metal3 ;
        RECT 269.505 12 270.165 12.66 ;
      LAYER Metal4 ;
        RECT 269.505 12 270.165 12.66 ;
    END
  END Q[18]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 272.385 12 273.045 12.66 ;
      LAYER Metal6 ;
        RECT 272.385 12 273.045 12.66 ;
      LAYER Metal3 ;
        RECT 272.385 12 273.045 12.66 ;
      LAYER Metal4 ;
        RECT 272.385 12 273.045 12.66 ;
    END
  END Q[19]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.94 12 26.6 12.66 ;
      LAYER Metal6 ;
        RECT 25.94 12 26.6 12.66 ;
      LAYER Metal3 ;
        RECT 25.94 12 26.6 12.66 ;
      LAYER Metal4 ;
        RECT 25.94 12 26.6 12.66 ;
    END
  END Q[1]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.845 12 292.505 12.66 ;
      LAYER Metal6 ;
        RECT 291.845 12 292.505 12.66 ;
      LAYER Metal3 ;
        RECT 291.845 12 292.505 12.66 ;
      LAYER Metal4 ;
        RECT 291.845 12 292.505 12.66 ;
    END
  END Q[20]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 294.725 12 295.385 12.66 ;
      LAYER Metal6 ;
        RECT 294.725 12 295.385 12.66 ;
      LAYER Metal3 ;
        RECT 294.725 12 295.385 12.66 ;
      LAYER Metal4 ;
        RECT 294.725 12 295.385 12.66 ;
    END
  END Q[21]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 313.125 12 313.785 12.66 ;
      LAYER Metal6 ;
        RECT 313.125 12 313.785 12.66 ;
      LAYER Metal3 ;
        RECT 313.125 12 313.785 12.66 ;
      LAYER Metal4 ;
        RECT 313.125 12 313.785 12.66 ;
    END
  END Q[22]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 316.005 12 316.665 12.66 ;
      LAYER Metal6 ;
        RECT 316.005 12 316.665 12.66 ;
      LAYER Metal3 ;
        RECT 316.005 12 316.665 12.66 ;
      LAYER Metal4 ;
        RECT 316.005 12 316.665 12.66 ;
    END
  END Q[23]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 335.465 12 336.125 12.66 ;
      LAYER Metal6 ;
        RECT 335.465 12 336.125 12.66 ;
      LAYER Metal3 ;
        RECT 335.465 12 336.125 12.66 ;
      LAYER Metal4 ;
        RECT 335.465 12 336.125 12.66 ;
    END
  END Q[24]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 338.345 12 339.005 12.66 ;
      LAYER Metal6 ;
        RECT 338.345 12 339.005 12.66 ;
      LAYER Metal3 ;
        RECT 338.345 12 339.005 12.66 ;
      LAYER Metal4 ;
        RECT 338.345 12 339.005 12.66 ;
    END
  END Q[25]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 356.745 12 357.405 12.66 ;
      LAYER Metal6 ;
        RECT 356.745 12 357.405 12.66 ;
      LAYER Metal3 ;
        RECT 356.745 12 357.405 12.66 ;
      LAYER Metal4 ;
        RECT 356.745 12 357.405 12.66 ;
    END
  END Q[26]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 359.625 12 360.285 12.66 ;
      LAYER Metal6 ;
        RECT 359.625 12 360.285 12.66 ;
      LAYER Metal3 ;
        RECT 359.625 12 360.285 12.66 ;
      LAYER Metal4 ;
        RECT 359.625 12 360.285 12.66 ;
    END
  END Q[27]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 379.085 12 379.745 12.66 ;
      LAYER Metal6 ;
        RECT 379.085 12 379.745 12.66 ;
      LAYER Metal3 ;
        RECT 379.085 12 379.745 12.66 ;
      LAYER Metal4 ;
        RECT 379.085 12 379.745 12.66 ;
    END
  END Q[28]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 381.965 12 382.625 12.66 ;
      LAYER Metal6 ;
        RECT 381.965 12 382.625 12.66 ;
      LAYER Metal3 ;
        RECT 381.965 12 382.625 12.66 ;
      LAYER Metal4 ;
        RECT 381.965 12 382.625 12.66 ;
    END
  END Q[29]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 44.34 12 45 12.66 ;
      LAYER Metal6 ;
        RECT 44.34 12 45 12.66 ;
      LAYER Metal3 ;
        RECT 44.34 12 45 12.66 ;
      LAYER Metal4 ;
        RECT 44.34 12 45 12.66 ;
    END
  END Q[2]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 400.365 12 401.025 12.66 ;
      LAYER Metal6 ;
        RECT 400.365 12 401.025 12.66 ;
      LAYER Metal3 ;
        RECT 400.365 12 401.025 12.66 ;
      LAYER Metal4 ;
        RECT 400.365 12 401.025 12.66 ;
    END
  END Q[30]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 403.245 12 403.905 12.66 ;
      LAYER Metal6 ;
        RECT 403.245 12 403.905 12.66 ;
      LAYER Metal3 ;
        RECT 403.245 12 403.905 12.66 ;
      LAYER Metal4 ;
        RECT 403.245 12 403.905 12.66 ;
    END
  END Q[31]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.22 12 47.88 12.66 ;
      LAYER Metal6 ;
        RECT 47.22 12 47.88 12.66 ;
      LAYER Metal3 ;
        RECT 47.22 12 47.88 12.66 ;
      LAYER Metal4 ;
        RECT 47.22 12 47.88 12.66 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 66.68 12 67.34 12.66 ;
      LAYER Metal6 ;
        RECT 66.68 12 67.34 12.66 ;
      LAYER Metal3 ;
        RECT 66.68 12 67.34 12.66 ;
      LAYER Metal4 ;
        RECT 66.68 12 67.34 12.66 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.56 12 70.22 12.66 ;
      LAYER Metal6 ;
        RECT 69.56 12 70.22 12.66 ;
      LAYER Metal3 ;
        RECT 69.56 12 70.22 12.66 ;
      LAYER Metal4 ;
        RECT 69.56 12 70.22 12.66 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 87.96 12 88.62 12.66 ;
      LAYER Metal6 ;
        RECT 87.96 12 88.62 12.66 ;
      LAYER Metal3 ;
        RECT 87.96 12 88.62 12.66 ;
      LAYER Metal4 ;
        RECT 87.96 12 88.62 12.66 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.84 12 91.5 12.66 ;
      LAYER Metal6 ;
        RECT 90.84 12 91.5 12.66 ;
      LAYER Metal3 ;
        RECT 90.84 12 91.5 12.66 ;
      LAYER Metal4 ;
        RECT 90.84 12 91.5 12.66 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.3 12 110.96 12.66 ;
      LAYER Metal6 ;
        RECT 110.3 12 110.96 12.66 ;
      LAYER Metal3 ;
        RECT 110.3 12 110.96 12.66 ;
      LAYER Metal4 ;
        RECT 110.3 12 110.96 12.66 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 113.18 12 113.84 12.66 ;
      LAYER Metal6 ;
        RECT 113.18 12 113.84 12.66 ;
      LAYER Metal3 ;
        RECT 113.18 12 113.84 12.66 ;
      LAYER Metal4 ;
        RECT 113.18 12 113.84 12.66 ;
    END
  END Q[9]
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 234.48 12 235.14 12.66 ;
      LAYER Metal6 ;
        RECT 234.48 12 235.14 12.66 ;
      LAYER Metal3 ;
        RECT 234.48 12 235.14 12.66 ;
      LAYER Metal4 ;
        RECT 234.48 12 235.14 12.66 ;
    END
  END WE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 109.215 426.965 114.215 ;
        RECT 0 0 426.965 5 ;
      LAYER Metal2 ;
        RECT 421.965 0 426.965 114.215 ;
        RECT 0 0 5 114.215 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 103.615 421.365 108.615 ;
        RECT 5.6 5.6 421.365 10.6 ;
      LAYER Metal2 ;
        RECT 416.365 5.6 421.365 108.615 ;
        RECT 5.6 5.6 10.6 108.615 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12 12 415.01 102.02 ;
    LAYER Metal2 ;
      RECT 12 12 415.01 102.02 ;
    LAYER Metal3 ;
      RECT 12 12 415.01 102.02 ;
    LAYER Metal4 ;
      RECT 12 12 415.01 102.02 ;
    LAYER Metal5 ;
      RECT 12 12 415.01 102.02 ;
    LAYER Metal6 ;
      RECT 12 12 415.01 102.02 ;
  END
END MEM1

MACRO MEM2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2 0 0 ;
  SIZE 423.015 BY 145.035 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 102.42 12.66 103.08 ;
      LAYER Metal6 ;
        RECT 12 102.42 12.66 103.08 ;
      LAYER Metal3 ;
        RECT 12 102.42 12.66 103.08 ;
      LAYER Metal4 ;
        RECT 12 102.42 12.66 103.08 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 96.3 12.66 96.96 ;
      LAYER Metal6 ;
        RECT 12 96.3 12.66 96.96 ;
      LAYER Metal3 ;
        RECT 12 96.3 12.66 96.96 ;
      LAYER Metal4 ;
        RECT 12 96.3 12.66 96.96 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 87.08 12.66 87.74 ;
      LAYER Metal6 ;
        RECT 12 87.08 12.66 87.74 ;
      LAYER Metal3 ;
        RECT 12 87.08 12.66 87.74 ;
      LAYER Metal4 ;
        RECT 12 87.08 12.66 87.74 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 84.06 12.66 84.72 ;
      LAYER Metal6 ;
        RECT 12 84.06 12.66 84.72 ;
      LAYER Metal3 ;
        RECT 12 84.06 12.66 84.72 ;
      LAYER Metal4 ;
        RECT 12 84.06 12.66 84.72 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 80.96 12.66 81.62 ;
      LAYER Metal6 ;
        RECT 12 80.96 12.66 81.62 ;
      LAYER Metal3 ;
        RECT 12 80.96 12.66 81.62 ;
      LAYER Metal4 ;
        RECT 12 80.96 12.66 81.62 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 74.84 12.66 75.5 ;
      LAYER Metal6 ;
        RECT 12 74.84 12.66 75.5 ;
      LAYER Metal3 ;
        RECT 12 74.84 12.66 75.5 ;
      LAYER Metal4 ;
        RECT 12 74.84 12.66 75.5 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 71.82 12.66 72.48 ;
      LAYER Metal6 ;
        RECT 12 71.82 12.66 72.48 ;
      LAYER Metal3 ;
        RECT 12 71.82 12.66 72.48 ;
      LAYER Metal4 ;
        RECT 12 71.82 12.66 72.48 ;
    END
  END A1[6]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 36.4 12.66 37.06 ;
      LAYER Metal6 ;
        RECT 12 36.4 12.66 37.06 ;
      LAYER Metal3 ;
        RECT 12 36.4 12.66 37.06 ;
      LAYER Metal4 ;
        RECT 12 36.4 12.66 37.06 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 42.52 12.66 43.18 ;
      LAYER Metal6 ;
        RECT 12 42.52 12.66 43.18 ;
      LAYER Metal3 ;
        RECT 12 42.52 12.66 43.18 ;
      LAYER Metal4 ;
        RECT 12 42.52 12.66 43.18 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 51.74 12.66 52.4 ;
      LAYER Metal6 ;
        RECT 12 51.74 12.66 52.4 ;
      LAYER Metal3 ;
        RECT 12 51.74 12.66 52.4 ;
      LAYER Metal4 ;
        RECT 12 51.74 12.66 52.4 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 54.76 12.66 55.42 ;
      LAYER Metal6 ;
        RECT 12 54.76 12.66 55.42 ;
      LAYER Metal3 ;
        RECT 12 54.76 12.66 55.42 ;
      LAYER Metal4 ;
        RECT 12 54.76 12.66 55.42 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 57.86 12.66 58.52 ;
      LAYER Metal6 ;
        RECT 12 57.86 12.66 58.52 ;
      LAYER Metal3 ;
        RECT 12 57.86 12.66 58.52 ;
      LAYER Metal4 ;
        RECT 12 57.86 12.66 58.52 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 63.98 12.66 64.64 ;
      LAYER Metal6 ;
        RECT 12 63.98 12.66 64.64 ;
      LAYER Metal3 ;
        RECT 12 63.98 12.66 64.64 ;
      LAYER Metal4 ;
        RECT 12 63.98 12.66 64.64 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 67 12.66 67.66 ;
      LAYER Metal6 ;
        RECT 12 67 12.66 67.66 ;
      LAYER Metal3 ;
        RECT 12 67 12.66 67.66 ;
      LAYER Metal4 ;
        RECT 12 67 12.66 67.66 ;
    END
  END A2[6]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 210.28 12 210.94 12.66 ;
      LAYER Metal6 ;
        RECT 210.28 12 210.94 12.66 ;
      LAYER Metal3 ;
        RECT 210.28 12 210.94 12.66 ;
      LAYER Metal4 ;
        RECT 210.28 12 210.94 12.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 196.36 12 197.02 12.66 ;
      LAYER Metal6 ;
        RECT 196.36 12 197.02 12.66 ;
      LAYER Metal3 ;
        RECT 196.36 12 197.02 12.66 ;
      LAYER Metal4 ;
        RECT 196.36 12 197.02 12.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 218.905 12 219.565 12.66 ;
      LAYER Metal6 ;
        RECT 218.905 12 219.565 12.66 ;
      LAYER Metal3 ;
        RECT 218.905 12 219.565 12.66 ;
      LAYER Metal4 ;
        RECT 218.905 12 219.565 12.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 187.735 12 188.395 12.66 ;
      LAYER Metal6 ;
        RECT 187.735 12 188.395 12.66 ;
      LAYER Metal3 ;
        RECT 187.735 12 188.395 12.66 ;
      LAYER Metal4 ;
        RECT 187.735 12 188.395 12.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 15.86 12 16.52 12.66 ;
      LAYER Metal6 ;
        RECT 15.86 12 16.52 12.66 ;
      LAYER Metal3 ;
        RECT 15.86 12 16.52 12.66 ;
      LAYER Metal4 ;
        RECT 15.86 12 16.52 12.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 122.26 12 122.92 12.66 ;
      LAYER Metal6 ;
        RECT 122.26 12 122.92 12.66 ;
      LAYER Metal3 ;
        RECT 122.26 12 122.92 12.66 ;
      LAYER Metal4 ;
        RECT 122.26 12 122.92 12.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 142.4 12 143.06 12.66 ;
      LAYER Metal6 ;
        RECT 142.4 12 143.06 12.66 ;
      LAYER Metal3 ;
        RECT 142.4 12 143.06 12.66 ;
      LAYER Metal4 ;
        RECT 142.4 12 143.06 12.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 143.54 12 144.2 12.66 ;
      LAYER Metal6 ;
        RECT 143.54 12 144.2 12.66 ;
      LAYER Metal3 ;
        RECT 143.54 12 144.2 12.66 ;
      LAYER Metal4 ;
        RECT 143.54 12 144.2 12.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 163.68 12 164.34 12.66 ;
      LAYER Metal6 ;
        RECT 163.68 12 164.34 12.66 ;
      LAYER Metal3 ;
        RECT 163.68 12 164.34 12.66 ;
      LAYER Metal4 ;
        RECT 163.68 12 164.34 12.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 164.82 12 165.48 12.66 ;
      LAYER Metal6 ;
        RECT 164.82 12 165.48 12.66 ;
      LAYER Metal3 ;
        RECT 164.82 12 165.48 12.66 ;
      LAYER Metal4 ;
        RECT 164.82 12 165.48 12.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 184.96 12 185.62 12.66 ;
      LAYER Metal6 ;
        RECT 184.96 12 185.62 12.66 ;
      LAYER Metal3 ;
        RECT 184.96 12 185.62 12.66 ;
      LAYER Metal4 ;
        RECT 184.96 12 185.62 12.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 221.68 12 222.34 12.66 ;
      LAYER Metal6 ;
        RECT 221.68 12 222.34 12.66 ;
      LAYER Metal3 ;
        RECT 221.68 12 222.34 12.66 ;
      LAYER Metal4 ;
        RECT 221.68 12 222.34 12.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 241.82 12 242.48 12.66 ;
      LAYER Metal6 ;
        RECT 241.82 12 242.48 12.66 ;
      LAYER Metal3 ;
        RECT 241.82 12 242.48 12.66 ;
      LAYER Metal4 ;
        RECT 241.82 12 242.48 12.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 242.96 12 243.62 12.66 ;
      LAYER Metal6 ;
        RECT 242.96 12 243.62 12.66 ;
      LAYER Metal3 ;
        RECT 242.96 12 243.62 12.66 ;
      LAYER Metal4 ;
        RECT 242.96 12 243.62 12.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 263.1 12 263.76 12.66 ;
      LAYER Metal6 ;
        RECT 263.1 12 263.76 12.66 ;
      LAYER Metal3 ;
        RECT 263.1 12 263.76 12.66 ;
      LAYER Metal4 ;
        RECT 263.1 12 263.76 12.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 36 12 36.66 12.66 ;
      LAYER Metal6 ;
        RECT 36 12 36.66 12.66 ;
      LAYER Metal3 ;
        RECT 36 12 36.66 12.66 ;
      LAYER Metal4 ;
        RECT 36 12 36.66 12.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 264.24 12 264.9 12.66 ;
      LAYER Metal6 ;
        RECT 264.24 12 264.9 12.66 ;
      LAYER Metal3 ;
        RECT 264.24 12 264.9 12.66 ;
      LAYER Metal4 ;
        RECT 264.24 12 264.9 12.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 284.38 12 285.04 12.66 ;
      LAYER Metal6 ;
        RECT 284.38 12 285.04 12.66 ;
      LAYER Metal3 ;
        RECT 284.38 12 285.04 12.66 ;
      LAYER Metal4 ;
        RECT 284.38 12 285.04 12.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 285.52 12 286.18 12.66 ;
      LAYER Metal6 ;
        RECT 285.52 12 286.18 12.66 ;
      LAYER Metal3 ;
        RECT 285.52 12 286.18 12.66 ;
      LAYER Metal4 ;
        RECT 285.52 12 286.18 12.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 305.66 12 306.32 12.66 ;
      LAYER Metal6 ;
        RECT 305.66 12 306.32 12.66 ;
      LAYER Metal3 ;
        RECT 305.66 12 306.32 12.66 ;
      LAYER Metal4 ;
        RECT 305.66 12 306.32 12.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 306.8 12 307.46 12.66 ;
      LAYER Metal6 ;
        RECT 306.8 12 307.46 12.66 ;
      LAYER Metal3 ;
        RECT 306.8 12 307.46 12.66 ;
      LAYER Metal4 ;
        RECT 306.8 12 307.46 12.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 326.94 12 327.6 12.66 ;
      LAYER Metal6 ;
        RECT 326.94 12 327.6 12.66 ;
      LAYER Metal3 ;
        RECT 326.94 12 327.6 12.66 ;
      LAYER Metal4 ;
        RECT 326.94 12 327.6 12.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 328.08 12 328.74 12.66 ;
      LAYER Metal6 ;
        RECT 328.08 12 328.74 12.66 ;
      LAYER Metal3 ;
        RECT 328.08 12 328.74 12.66 ;
      LAYER Metal4 ;
        RECT 328.08 12 328.74 12.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 348.22 12 348.88 12.66 ;
      LAYER Metal6 ;
        RECT 348.22 12 348.88 12.66 ;
      LAYER Metal3 ;
        RECT 348.22 12 348.88 12.66 ;
      LAYER Metal4 ;
        RECT 348.22 12 348.88 12.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 349.36 12 350.02 12.66 ;
      LAYER Metal6 ;
        RECT 349.36 12 350.02 12.66 ;
      LAYER Metal3 ;
        RECT 349.36 12 350.02 12.66 ;
      LAYER Metal4 ;
        RECT 349.36 12 350.02 12.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 369.5 12 370.16 12.66 ;
      LAYER Metal6 ;
        RECT 369.5 12 370.16 12.66 ;
      LAYER Metal3 ;
        RECT 369.5 12 370.16 12.66 ;
      LAYER Metal4 ;
        RECT 369.5 12 370.16 12.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 37.14 12 37.8 12.66 ;
      LAYER Metal6 ;
        RECT 37.14 12 37.8 12.66 ;
      LAYER Metal3 ;
        RECT 37.14 12 37.8 12.66 ;
      LAYER Metal4 ;
        RECT 37.14 12 37.8 12.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 370.64 12 371.3 12.66 ;
      LAYER Metal6 ;
        RECT 370.64 12 371.3 12.66 ;
      LAYER Metal3 ;
        RECT 370.64 12 371.3 12.66 ;
      LAYER Metal4 ;
        RECT 370.64 12 371.3 12.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 390.78 12 391.44 12.66 ;
      LAYER Metal6 ;
        RECT 390.78 12 391.44 12.66 ;
      LAYER Metal3 ;
        RECT 390.78 12 391.44 12.66 ;
      LAYER Metal4 ;
        RECT 390.78 12 391.44 12.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 57.28 12 57.94 12.66 ;
      LAYER Metal6 ;
        RECT 57.28 12 57.94 12.66 ;
      LAYER Metal3 ;
        RECT 57.28 12 57.94 12.66 ;
      LAYER Metal4 ;
        RECT 57.28 12 57.94 12.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 58.42 12 59.08 12.66 ;
      LAYER Metal6 ;
        RECT 58.42 12 59.08 12.66 ;
      LAYER Metal3 ;
        RECT 58.42 12 59.08 12.66 ;
      LAYER Metal4 ;
        RECT 58.42 12 59.08 12.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 78.56 12 79.22 12.66 ;
      LAYER Metal6 ;
        RECT 78.56 12 79.22 12.66 ;
      LAYER Metal3 ;
        RECT 78.56 12 79.22 12.66 ;
      LAYER Metal4 ;
        RECT 78.56 12 79.22 12.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 79.7 12 80.36 12.66 ;
      LAYER Metal6 ;
        RECT 79.7 12 80.36 12.66 ;
      LAYER Metal3 ;
        RECT 79.7 12 80.36 12.66 ;
      LAYER Metal4 ;
        RECT 79.7 12 80.36 12.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 99.84 12 100.5 12.66 ;
      LAYER Metal6 ;
        RECT 99.84 12 100.5 12.66 ;
      LAYER Metal3 ;
        RECT 99.84 12 100.5 12.66 ;
      LAYER Metal4 ;
        RECT 99.84 12 100.5 12.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 100.98 12 101.64 12.66 ;
      LAYER Metal6 ;
        RECT 100.98 12 101.64 12.66 ;
      LAYER Metal3 ;
        RECT 100.98 12 101.64 12.66 ;
      LAYER Metal4 ;
        RECT 100.98 12 101.64 12.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 121.12 12 121.78 12.66 ;
      LAYER Metal6 ;
        RECT 121.12 12 121.78 12.66 ;
      LAYER Metal3 ;
        RECT 121.12 12 121.78 12.66 ;
      LAYER Metal4 ;
        RECT 121.12 12 121.78 12.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.36 12 26.02 12.66 ;
      LAYER Metal6 ;
        RECT 25.36 12 26.02 12.66 ;
      LAYER Metal3 ;
        RECT 25.36 12 26.02 12.66 ;
      LAYER Metal4 ;
        RECT 25.36 12 26.02 12.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.76 12 132.42 12.66 ;
      LAYER Metal6 ;
        RECT 131.76 12 132.42 12.66 ;
      LAYER Metal3 ;
        RECT 131.76 12 132.42 12.66 ;
      LAYER Metal4 ;
        RECT 131.76 12 132.42 12.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 132.9 12 133.56 12.66 ;
      LAYER Metal6 ;
        RECT 132.9 12 133.56 12.66 ;
      LAYER Metal3 ;
        RECT 132.9 12 133.56 12.66 ;
      LAYER Metal4 ;
        RECT 132.9 12 133.56 12.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.04 12 153.7 12.66 ;
      LAYER Metal6 ;
        RECT 153.04 12 153.7 12.66 ;
      LAYER Metal3 ;
        RECT 153.04 12 153.7 12.66 ;
      LAYER Metal4 ;
        RECT 153.04 12 153.7 12.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 154.18 12 154.84 12.66 ;
      LAYER Metal6 ;
        RECT 154.18 12 154.84 12.66 ;
      LAYER Metal3 ;
        RECT 154.18 12 154.84 12.66 ;
      LAYER Metal4 ;
        RECT 154.18 12 154.84 12.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 174.32 12 174.98 12.66 ;
      LAYER Metal6 ;
        RECT 174.32 12 174.98 12.66 ;
      LAYER Metal3 ;
        RECT 174.32 12 174.98 12.66 ;
      LAYER Metal4 ;
        RECT 174.32 12 174.98 12.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.46 12 176.12 12.66 ;
      LAYER Metal6 ;
        RECT 175.46 12 176.12 12.66 ;
      LAYER Metal3 ;
        RECT 175.46 12 176.12 12.66 ;
      LAYER Metal4 ;
        RECT 175.46 12 176.12 12.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 231.18 12 231.84 12.66 ;
      LAYER Metal6 ;
        RECT 231.18 12 231.84 12.66 ;
      LAYER Metal3 ;
        RECT 231.18 12 231.84 12.66 ;
      LAYER Metal4 ;
        RECT 231.18 12 231.84 12.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 232.32 12 232.98 12.66 ;
      LAYER Metal6 ;
        RECT 232.32 12 232.98 12.66 ;
      LAYER Metal3 ;
        RECT 232.32 12 232.98 12.66 ;
      LAYER Metal4 ;
        RECT 232.32 12 232.98 12.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 252.46 12 253.12 12.66 ;
      LAYER Metal6 ;
        RECT 252.46 12 253.12 12.66 ;
      LAYER Metal3 ;
        RECT 252.46 12 253.12 12.66 ;
      LAYER Metal4 ;
        RECT 252.46 12 253.12 12.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 253.6 12 254.26 12.66 ;
      LAYER Metal6 ;
        RECT 253.6 12 254.26 12.66 ;
      LAYER Metal3 ;
        RECT 253.6 12 254.26 12.66 ;
      LAYER Metal4 ;
        RECT 253.6 12 254.26 12.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 26.5 12 27.16 12.66 ;
      LAYER Metal6 ;
        RECT 26.5 12 27.16 12.66 ;
      LAYER Metal3 ;
        RECT 26.5 12 27.16 12.66 ;
      LAYER Metal4 ;
        RECT 26.5 12 27.16 12.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 273.74 12 274.4 12.66 ;
      LAYER Metal6 ;
        RECT 273.74 12 274.4 12.66 ;
      LAYER Metal3 ;
        RECT 273.74 12 274.4 12.66 ;
      LAYER Metal4 ;
        RECT 273.74 12 274.4 12.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 274.88 12 275.54 12.66 ;
      LAYER Metal6 ;
        RECT 274.88 12 275.54 12.66 ;
      LAYER Metal3 ;
        RECT 274.88 12 275.54 12.66 ;
      LAYER Metal4 ;
        RECT 274.88 12 275.54 12.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 295.02 12 295.68 12.66 ;
      LAYER Metal6 ;
        RECT 295.02 12 295.68 12.66 ;
      LAYER Metal3 ;
        RECT 295.02 12 295.68 12.66 ;
      LAYER Metal4 ;
        RECT 295.02 12 295.68 12.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 296.16 12 296.82 12.66 ;
      LAYER Metal6 ;
        RECT 296.16 12 296.82 12.66 ;
      LAYER Metal3 ;
        RECT 296.16 12 296.82 12.66 ;
      LAYER Metal4 ;
        RECT 296.16 12 296.82 12.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 316.3 12 316.96 12.66 ;
      LAYER Metal6 ;
        RECT 316.3 12 316.96 12.66 ;
      LAYER Metal3 ;
        RECT 316.3 12 316.96 12.66 ;
      LAYER Metal4 ;
        RECT 316.3 12 316.96 12.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 317.44 12 318.1 12.66 ;
      LAYER Metal6 ;
        RECT 317.44 12 318.1 12.66 ;
      LAYER Metal3 ;
        RECT 317.44 12 318.1 12.66 ;
      LAYER Metal4 ;
        RECT 317.44 12 318.1 12.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 337.58 12 338.24 12.66 ;
      LAYER Metal6 ;
        RECT 337.58 12 338.24 12.66 ;
      LAYER Metal3 ;
        RECT 337.58 12 338.24 12.66 ;
      LAYER Metal4 ;
        RECT 337.58 12 338.24 12.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 338.72 12 339.38 12.66 ;
      LAYER Metal6 ;
        RECT 338.72 12 339.38 12.66 ;
      LAYER Metal3 ;
        RECT 338.72 12 339.38 12.66 ;
      LAYER Metal4 ;
        RECT 338.72 12 339.38 12.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 358.86 12 359.52 12.66 ;
      LAYER Metal6 ;
        RECT 358.86 12 359.52 12.66 ;
      LAYER Metal3 ;
        RECT 358.86 12 359.52 12.66 ;
      LAYER Metal4 ;
        RECT 358.86 12 359.52 12.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 360 12 360.66 12.66 ;
      LAYER Metal6 ;
        RECT 360 12 360.66 12.66 ;
      LAYER Metal3 ;
        RECT 360 12 360.66 12.66 ;
      LAYER Metal4 ;
        RECT 360 12 360.66 12.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 46.64 12 47.3 12.66 ;
      LAYER Metal6 ;
        RECT 46.64 12 47.3 12.66 ;
      LAYER Metal3 ;
        RECT 46.64 12 47.3 12.66 ;
      LAYER Metal4 ;
        RECT 46.64 12 47.3 12.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 380.14 12 380.8 12.66 ;
      LAYER Metal6 ;
        RECT 380.14 12 380.8 12.66 ;
      LAYER Metal3 ;
        RECT 380.14 12 380.8 12.66 ;
      LAYER Metal4 ;
        RECT 380.14 12 380.8 12.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 381.28 12 381.94 12.66 ;
      LAYER Metal6 ;
        RECT 381.28 12 381.94 12.66 ;
      LAYER Metal3 ;
        RECT 381.28 12 381.94 12.66 ;
      LAYER Metal4 ;
        RECT 381.28 12 381.94 12.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.78 12 48.44 12.66 ;
      LAYER Metal6 ;
        RECT 47.78 12 48.44 12.66 ;
      LAYER Metal3 ;
        RECT 47.78 12 48.44 12.66 ;
      LAYER Metal4 ;
        RECT 47.78 12 48.44 12.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 67.92 12 68.58 12.66 ;
      LAYER Metal6 ;
        RECT 67.92 12 68.58 12.66 ;
      LAYER Metal3 ;
        RECT 67.92 12 68.58 12.66 ;
      LAYER Metal4 ;
        RECT 67.92 12 68.58 12.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.06 12 69.72 12.66 ;
      LAYER Metal6 ;
        RECT 69.06 12 69.72 12.66 ;
      LAYER Metal3 ;
        RECT 69.06 12 69.72 12.66 ;
      LAYER Metal4 ;
        RECT 69.06 12 69.72 12.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 89.2 12 89.86 12.66 ;
      LAYER Metal6 ;
        RECT 89.2 12 89.86 12.66 ;
      LAYER Metal3 ;
        RECT 89.2 12 89.86 12.66 ;
      LAYER Metal4 ;
        RECT 89.2 12 89.86 12.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.34 12 91 12.66 ;
      LAYER Metal6 ;
        RECT 90.34 12 91 12.66 ;
      LAYER Metal3 ;
        RECT 90.34 12 91 12.66 ;
      LAYER Metal4 ;
        RECT 90.34 12 91 12.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.48 12 111.14 12.66 ;
      LAYER Metal6 ;
        RECT 110.48 12 111.14 12.66 ;
      LAYER Metal3 ;
        RECT 110.48 12 111.14 12.66 ;
      LAYER Metal4 ;
        RECT 110.48 12 111.14 12.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 111.62 12 112.28 12.66 ;
      LAYER Metal6 ;
        RECT 111.62 12 112.28 12.66 ;
      LAYER Metal3 ;
        RECT 111.62 12 112.28 12.66 ;
      LAYER Metal4 ;
        RECT 111.62 12 112.28 12.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 18.28 12 18.94 12.66 ;
      LAYER Metal6 ;
        RECT 18.28 12 18.94 12.66 ;
      LAYER Metal3 ;
        RECT 18.28 12 18.94 12.66 ;
      LAYER Metal4 ;
        RECT 18.28 12 18.94 12.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 125.56 12 126.22 12.66 ;
      LAYER Metal6 ;
        RECT 125.56 12 126.22 12.66 ;
      LAYER Metal3 ;
        RECT 125.56 12 126.22 12.66 ;
      LAYER Metal4 ;
        RECT 125.56 12 126.22 12.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 139.1 12 139.76 12.66 ;
      LAYER Metal6 ;
        RECT 139.1 12 139.76 12.66 ;
      LAYER Metal3 ;
        RECT 139.1 12 139.76 12.66 ;
      LAYER Metal4 ;
        RECT 139.1 12 139.76 12.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 146.84 12 147.5 12.66 ;
      LAYER Metal6 ;
        RECT 146.84 12 147.5 12.66 ;
      LAYER Metal3 ;
        RECT 146.84 12 147.5 12.66 ;
      LAYER Metal4 ;
        RECT 146.84 12 147.5 12.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 160.38 12 161.04 12.66 ;
      LAYER Metal6 ;
        RECT 160.38 12 161.04 12.66 ;
      LAYER Metal3 ;
        RECT 160.38 12 161.04 12.66 ;
      LAYER Metal4 ;
        RECT 160.38 12 161.04 12.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 168.12 12 168.78 12.66 ;
      LAYER Metal6 ;
        RECT 168.12 12 168.78 12.66 ;
      LAYER Metal3 ;
        RECT 168.12 12 168.78 12.66 ;
      LAYER Metal4 ;
        RECT 168.12 12 168.78 12.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 181.66 12 182.32 12.66 ;
      LAYER Metal6 ;
        RECT 181.66 12 182.32 12.66 ;
      LAYER Metal3 ;
        RECT 181.66 12 182.32 12.66 ;
      LAYER Metal4 ;
        RECT 181.66 12 182.32 12.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 224.98 12 225.64 12.66 ;
      LAYER Metal6 ;
        RECT 224.98 12 225.64 12.66 ;
      LAYER Metal3 ;
        RECT 224.98 12 225.64 12.66 ;
      LAYER Metal4 ;
        RECT 224.98 12 225.64 12.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 238.52 12 239.18 12.66 ;
      LAYER Metal6 ;
        RECT 238.52 12 239.18 12.66 ;
      LAYER Metal3 ;
        RECT 238.52 12 239.18 12.66 ;
      LAYER Metal4 ;
        RECT 238.52 12 239.18 12.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 246.26 12 246.92 12.66 ;
      LAYER Metal6 ;
        RECT 246.26 12 246.92 12.66 ;
      LAYER Metal3 ;
        RECT 246.26 12 246.92 12.66 ;
      LAYER Metal4 ;
        RECT 246.26 12 246.92 12.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 259.8 12 260.46 12.66 ;
      LAYER Metal6 ;
        RECT 259.8 12 260.46 12.66 ;
      LAYER Metal3 ;
        RECT 259.8 12 260.46 12.66 ;
      LAYER Metal4 ;
        RECT 259.8 12 260.46 12.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 32.7 12 33.36 12.66 ;
      LAYER Metal6 ;
        RECT 32.7 12 33.36 12.66 ;
      LAYER Metal3 ;
        RECT 32.7 12 33.36 12.66 ;
      LAYER Metal4 ;
        RECT 32.7 12 33.36 12.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 267.54 12 268.2 12.66 ;
      LAYER Metal6 ;
        RECT 267.54 12 268.2 12.66 ;
      LAYER Metal3 ;
        RECT 267.54 12 268.2 12.66 ;
      LAYER Metal4 ;
        RECT 267.54 12 268.2 12.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 281.08 12 281.74 12.66 ;
      LAYER Metal6 ;
        RECT 281.08 12 281.74 12.66 ;
      LAYER Metal3 ;
        RECT 281.08 12 281.74 12.66 ;
      LAYER Metal4 ;
        RECT 281.08 12 281.74 12.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 288.82 12 289.48 12.66 ;
      LAYER Metal6 ;
        RECT 288.82 12 289.48 12.66 ;
      LAYER Metal3 ;
        RECT 288.82 12 289.48 12.66 ;
      LAYER Metal4 ;
        RECT 288.82 12 289.48 12.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 302.36 12 303.02 12.66 ;
      LAYER Metal6 ;
        RECT 302.36 12 303.02 12.66 ;
      LAYER Metal3 ;
        RECT 302.36 12 303.02 12.66 ;
      LAYER Metal4 ;
        RECT 302.36 12 303.02 12.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 310.1 12 310.76 12.66 ;
      LAYER Metal6 ;
        RECT 310.1 12 310.76 12.66 ;
      LAYER Metal3 ;
        RECT 310.1 12 310.76 12.66 ;
      LAYER Metal4 ;
        RECT 310.1 12 310.76 12.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 323.64 12 324.3 12.66 ;
      LAYER Metal6 ;
        RECT 323.64 12 324.3 12.66 ;
      LAYER Metal3 ;
        RECT 323.64 12 324.3 12.66 ;
      LAYER Metal4 ;
        RECT 323.64 12 324.3 12.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 331.38 12 332.04 12.66 ;
      LAYER Metal6 ;
        RECT 331.38 12 332.04 12.66 ;
      LAYER Metal3 ;
        RECT 331.38 12 332.04 12.66 ;
      LAYER Metal4 ;
        RECT 331.38 12 332.04 12.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 344.92 12 345.58 12.66 ;
      LAYER Metal6 ;
        RECT 344.92 12 345.58 12.66 ;
      LAYER Metal3 ;
        RECT 344.92 12 345.58 12.66 ;
      LAYER Metal4 ;
        RECT 344.92 12 345.58 12.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 352.66 12 353.32 12.66 ;
      LAYER Metal6 ;
        RECT 352.66 12 353.32 12.66 ;
      LAYER Metal3 ;
        RECT 352.66 12 353.32 12.66 ;
      LAYER Metal4 ;
        RECT 352.66 12 353.32 12.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 366.2 12 366.86 12.66 ;
      LAYER Metal6 ;
        RECT 366.2 12 366.86 12.66 ;
      LAYER Metal3 ;
        RECT 366.2 12 366.86 12.66 ;
      LAYER Metal4 ;
        RECT 366.2 12 366.86 12.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 40.44 12 41.1 12.66 ;
      LAYER Metal6 ;
        RECT 40.44 12 41.1 12.66 ;
      LAYER Metal3 ;
        RECT 40.44 12 41.1 12.66 ;
      LAYER Metal4 ;
        RECT 40.44 12 41.1 12.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 373.94 12 374.6 12.66 ;
      LAYER Metal6 ;
        RECT 373.94 12 374.6 12.66 ;
      LAYER Metal3 ;
        RECT 373.94 12 374.6 12.66 ;
      LAYER Metal4 ;
        RECT 373.94 12 374.6 12.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 388.36 12 389.02 12.66 ;
      LAYER Metal6 ;
        RECT 388.36 12 389.02 12.66 ;
      LAYER Metal3 ;
        RECT 388.36 12 389.02 12.66 ;
      LAYER Metal4 ;
        RECT 388.36 12 389.02 12.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 53.98 12 54.64 12.66 ;
      LAYER Metal6 ;
        RECT 53.98 12 54.64 12.66 ;
      LAYER Metal3 ;
        RECT 53.98 12 54.64 12.66 ;
      LAYER Metal4 ;
        RECT 53.98 12 54.64 12.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 61.72 12 62.38 12.66 ;
      LAYER Metal6 ;
        RECT 61.72 12 62.38 12.66 ;
      LAYER Metal3 ;
        RECT 61.72 12 62.38 12.66 ;
      LAYER Metal4 ;
        RECT 61.72 12 62.38 12.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 75.26 12 75.92 12.66 ;
      LAYER Metal6 ;
        RECT 75.26 12 75.92 12.66 ;
      LAYER Metal3 ;
        RECT 75.26 12 75.92 12.66 ;
      LAYER Metal4 ;
        RECT 75.26 12 75.92 12.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 83 12 83.66 12.66 ;
      LAYER Metal6 ;
        RECT 83 12 83.66 12.66 ;
      LAYER Metal3 ;
        RECT 83 12 83.66 12.66 ;
      LAYER Metal4 ;
        RECT 83 12 83.66 12.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 96.54 12 97.2 12.66 ;
      LAYER Metal6 ;
        RECT 96.54 12 97.2 12.66 ;
      LAYER Metal3 ;
        RECT 96.54 12 97.2 12.66 ;
      LAYER Metal4 ;
        RECT 96.54 12 97.2 12.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 104.28 12 104.94 12.66 ;
      LAYER Metal6 ;
        RECT 104.28 12 104.94 12.66 ;
      LAYER Metal3 ;
        RECT 104.28 12 104.94 12.66 ;
      LAYER Metal4 ;
        RECT 104.28 12 104.94 12.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 117.82 12 118.48 12.66 ;
      LAYER Metal6 ;
        RECT 117.82 12 118.48 12.66 ;
      LAYER Metal3 ;
        RECT 117.82 12 118.48 12.66 ;
      LAYER Metal4 ;
        RECT 117.82 12 118.48 12.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 22.06 12 22.72 12.66 ;
      LAYER Metal6 ;
        RECT 22.06 12 22.72 12.66 ;
      LAYER Metal3 ;
        RECT 22.06 12 22.72 12.66 ;
      LAYER Metal4 ;
        RECT 22.06 12 22.72 12.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 128.46 12 129.12 12.66 ;
      LAYER Metal6 ;
        RECT 128.46 12 129.12 12.66 ;
      LAYER Metal3 ;
        RECT 128.46 12 129.12 12.66 ;
      LAYER Metal4 ;
        RECT 128.46 12 129.12 12.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 136.2 12 136.86 12.66 ;
      LAYER Metal6 ;
        RECT 136.2 12 136.86 12.66 ;
      LAYER Metal3 ;
        RECT 136.2 12 136.86 12.66 ;
      LAYER Metal4 ;
        RECT 136.2 12 136.86 12.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 149.74 12 150.4 12.66 ;
      LAYER Metal6 ;
        RECT 149.74 12 150.4 12.66 ;
      LAYER Metal3 ;
        RECT 149.74 12 150.4 12.66 ;
      LAYER Metal4 ;
        RECT 149.74 12 150.4 12.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 157.48 12 158.14 12.66 ;
      LAYER Metal6 ;
        RECT 157.48 12 158.14 12.66 ;
      LAYER Metal3 ;
        RECT 157.48 12 158.14 12.66 ;
      LAYER Metal4 ;
        RECT 157.48 12 158.14 12.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 171.02 12 171.68 12.66 ;
      LAYER Metal6 ;
        RECT 171.02 12 171.68 12.66 ;
      LAYER Metal3 ;
        RECT 171.02 12 171.68 12.66 ;
      LAYER Metal4 ;
        RECT 171.02 12 171.68 12.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.76 12 179.42 12.66 ;
      LAYER Metal6 ;
        RECT 178.76 12 179.42 12.66 ;
      LAYER Metal3 ;
        RECT 178.76 12 179.42 12.66 ;
      LAYER Metal4 ;
        RECT 178.76 12 179.42 12.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 227.88 12 228.54 12.66 ;
      LAYER Metal6 ;
        RECT 227.88 12 228.54 12.66 ;
      LAYER Metal3 ;
        RECT 227.88 12 228.54 12.66 ;
      LAYER Metal4 ;
        RECT 227.88 12 228.54 12.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 235.62 12 236.28 12.66 ;
      LAYER Metal6 ;
        RECT 235.62 12 236.28 12.66 ;
      LAYER Metal3 ;
        RECT 235.62 12 236.28 12.66 ;
      LAYER Metal4 ;
        RECT 235.62 12 236.28 12.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 249.16 12 249.82 12.66 ;
      LAYER Metal6 ;
        RECT 249.16 12 249.82 12.66 ;
      LAYER Metal3 ;
        RECT 249.16 12 249.82 12.66 ;
      LAYER Metal4 ;
        RECT 249.16 12 249.82 12.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 256.9 12 257.56 12.66 ;
      LAYER Metal6 ;
        RECT 256.9 12 257.56 12.66 ;
      LAYER Metal3 ;
        RECT 256.9 12 257.56 12.66 ;
      LAYER Metal4 ;
        RECT 256.9 12 257.56 12.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 29.8 12 30.46 12.66 ;
      LAYER Metal6 ;
        RECT 29.8 12 30.46 12.66 ;
      LAYER Metal3 ;
        RECT 29.8 12 30.46 12.66 ;
      LAYER Metal4 ;
        RECT 29.8 12 30.46 12.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 270.44 12 271.1 12.66 ;
      LAYER Metal6 ;
        RECT 270.44 12 271.1 12.66 ;
      LAYER Metal3 ;
        RECT 270.44 12 271.1 12.66 ;
      LAYER Metal4 ;
        RECT 270.44 12 271.1 12.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 278.18 12 278.84 12.66 ;
      LAYER Metal6 ;
        RECT 278.18 12 278.84 12.66 ;
      LAYER Metal3 ;
        RECT 278.18 12 278.84 12.66 ;
      LAYER Metal4 ;
        RECT 278.18 12 278.84 12.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.72 12 292.38 12.66 ;
      LAYER Metal6 ;
        RECT 291.72 12 292.38 12.66 ;
      LAYER Metal3 ;
        RECT 291.72 12 292.38 12.66 ;
      LAYER Metal4 ;
        RECT 291.72 12 292.38 12.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 299.46 12 300.12 12.66 ;
      LAYER Metal6 ;
        RECT 299.46 12 300.12 12.66 ;
      LAYER Metal3 ;
        RECT 299.46 12 300.12 12.66 ;
      LAYER Metal4 ;
        RECT 299.46 12 300.12 12.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 313 12 313.66 12.66 ;
      LAYER Metal6 ;
        RECT 313 12 313.66 12.66 ;
      LAYER Metal3 ;
        RECT 313 12 313.66 12.66 ;
      LAYER Metal4 ;
        RECT 313 12 313.66 12.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 320.74 12 321.4 12.66 ;
      LAYER Metal6 ;
        RECT 320.74 12 321.4 12.66 ;
      LAYER Metal3 ;
        RECT 320.74 12 321.4 12.66 ;
      LAYER Metal4 ;
        RECT 320.74 12 321.4 12.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 334.28 12 334.94 12.66 ;
      LAYER Metal6 ;
        RECT 334.28 12 334.94 12.66 ;
      LAYER Metal3 ;
        RECT 334.28 12 334.94 12.66 ;
      LAYER Metal4 ;
        RECT 334.28 12 334.94 12.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 342.02 12 342.68 12.66 ;
      LAYER Metal6 ;
        RECT 342.02 12 342.68 12.66 ;
      LAYER Metal3 ;
        RECT 342.02 12 342.68 12.66 ;
      LAYER Metal4 ;
        RECT 342.02 12 342.68 12.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 355.56 12 356.22 12.66 ;
      LAYER Metal6 ;
        RECT 355.56 12 356.22 12.66 ;
      LAYER Metal3 ;
        RECT 355.56 12 356.22 12.66 ;
      LAYER Metal4 ;
        RECT 355.56 12 356.22 12.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 363.3 12 363.96 12.66 ;
      LAYER Metal6 ;
        RECT 363.3 12 363.96 12.66 ;
      LAYER Metal3 ;
        RECT 363.3 12 363.96 12.66 ;
      LAYER Metal4 ;
        RECT 363.3 12 363.96 12.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 43.34 12 44 12.66 ;
      LAYER Metal6 ;
        RECT 43.34 12 44 12.66 ;
      LAYER Metal3 ;
        RECT 43.34 12 44 12.66 ;
      LAYER Metal4 ;
        RECT 43.34 12 44 12.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.84 12 377.5 12.66 ;
      LAYER Metal6 ;
        RECT 376.84 12 377.5 12.66 ;
      LAYER Metal3 ;
        RECT 376.84 12 377.5 12.66 ;
      LAYER Metal4 ;
        RECT 376.84 12 377.5 12.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.58 12 385.24 12.66 ;
      LAYER Metal6 ;
        RECT 384.58 12 385.24 12.66 ;
      LAYER Metal3 ;
        RECT 384.58 12 385.24 12.66 ;
      LAYER Metal4 ;
        RECT 384.58 12 385.24 12.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 51.08 12 51.74 12.66 ;
      LAYER Metal6 ;
        RECT 51.08 12 51.74 12.66 ;
      LAYER Metal3 ;
        RECT 51.08 12 51.74 12.66 ;
      LAYER Metal4 ;
        RECT 51.08 12 51.74 12.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.62 12 65.28 12.66 ;
      LAYER Metal6 ;
        RECT 64.62 12 65.28 12.66 ;
      LAYER Metal3 ;
        RECT 64.62 12 65.28 12.66 ;
      LAYER Metal4 ;
        RECT 64.62 12 65.28 12.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.36 12 73.02 12.66 ;
      LAYER Metal6 ;
        RECT 72.36 12 73.02 12.66 ;
      LAYER Metal3 ;
        RECT 72.36 12 73.02 12.66 ;
      LAYER Metal4 ;
        RECT 72.36 12 73.02 12.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.9 12 86.56 12.66 ;
      LAYER Metal6 ;
        RECT 85.9 12 86.56 12.66 ;
      LAYER Metal3 ;
        RECT 85.9 12 86.56 12.66 ;
      LAYER Metal4 ;
        RECT 85.9 12 86.56 12.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.64 12 94.3 12.66 ;
      LAYER Metal6 ;
        RECT 93.64 12 94.3 12.66 ;
      LAYER Metal3 ;
        RECT 93.64 12 94.3 12.66 ;
      LAYER Metal4 ;
        RECT 93.64 12 94.3 12.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.18 12 107.84 12.66 ;
      LAYER Metal6 ;
        RECT 107.18 12 107.84 12.66 ;
      LAYER Metal3 ;
        RECT 107.18 12 107.84 12.66 ;
      LAYER Metal4 ;
        RECT 107.18 12 107.84 12.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 114.92 12 115.58 12.66 ;
      LAYER Metal6 ;
        RECT 114.92 12 115.58 12.66 ;
      LAYER Metal3 ;
        RECT 114.92 12 115.58 12.66 ;
      LAYER Metal4 ;
        RECT 114.92 12 115.58 12.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 212.68 12 213.34 12.66 ;
      LAYER Metal6 ;
        RECT 212.68 12 213.34 12.66 ;
      LAYER Metal3 ;
        RECT 212.68 12 213.34 12.66 ;
      LAYER Metal4 ;
        RECT 212.68 12 213.34 12.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 193.96 12 194.62 12.66 ;
      LAYER Metal6 ;
        RECT 193.96 12 194.62 12.66 ;
      LAYER Metal3 ;
        RECT 193.96 12 194.62 12.66 ;
      LAYER Metal4 ;
        RECT 193.96 12 194.62 12.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 140.035 423.015 145.035 ;
        RECT 0 0 423.015 5 ;
      LAYER Metal2 ;
        RECT 418.015 0 423.015 145.035 ;
        RECT 0 0 5 145.035 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 134.435 417.415 139.435 ;
        RECT 5.6 5.6 417.415 10.6 ;
      LAYER Metal2 ;
        RECT 412.415 5.6 417.415 139.435 ;
        RECT 5.6 5.6 10.6 139.435 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal2 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal3 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal4 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal5 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal6 ;
      RECT 12 12 411.02 132.965 ;
  END
END MEM2

END LIBRARY
